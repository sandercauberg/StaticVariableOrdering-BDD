//# 35 inputs
//# 320 outputs
//# 1728 D-type flipflops
//# 3861 inverters
//# 12204 gates (4032 ANDs + 7020 NANDs + 1152 ORs + 0 NORs)

module dff (CK,Q,D);
input CK,D;
output Q;

  wire NM,NCK;
  trireg NQ,M;

  nmos N7 (M,D,NCK);
  not P3 (NM,M);
  nmos N9 (NQ,NM,CK);
  not P5 (Q,NQ);
  not P1 (NCK,CK);

endmodule

module s35932(GND,VDD,CK,CRC_OUT_1_0,CRC_OUT_1_1,CRC_OUT_1_10,CRC_OUT_1_11,
  CRC_OUT_1_12,CRC_OUT_1_13,CRC_OUT_1_14,CRC_OUT_1_15,CRC_OUT_1_16,CRC_OUT_1_17,
  CRC_OUT_1_18,CRC_OUT_1_19,CRC_OUT_1_2,CRC_OUT_1_20,CRC_OUT_1_21,CRC_OUT_1_22,
  CRC_OUT_1_23,CRC_OUT_1_24,CRC_OUT_1_25,CRC_OUT_1_26,CRC_OUT_1_27,
  CRC_OUT_1_28,CRC_OUT_1_29,CRC_OUT_1_3,CRC_OUT_1_30,CRC_OUT_1_31,CRC_OUT_1_4,
  CRC_OUT_1_5,CRC_OUT_1_6,CRC_OUT_1_7,CRC_OUT_1_8,CRC_OUT_1_9,CRC_OUT_2_0,
  CRC_OUT_2_1,CRC_OUT_2_10,CRC_OUT_2_11,CRC_OUT_2_12,CRC_OUT_2_13,CRC_OUT_2_14,
  CRC_OUT_2_15,CRC_OUT_2_16,CRC_OUT_2_17,CRC_OUT_2_18,CRC_OUT_2_19,CRC_OUT_2_2,
  CRC_OUT_2_20,CRC_OUT_2_21,CRC_OUT_2_22,CRC_OUT_2_23,CRC_OUT_2_24,
  CRC_OUT_2_25,CRC_OUT_2_26,CRC_OUT_2_27,CRC_OUT_2_28,CRC_OUT_2_29,CRC_OUT_2_3,
  CRC_OUT_2_30,CRC_OUT_2_31,CRC_OUT_2_4,CRC_OUT_2_5,CRC_OUT_2_6,CRC_OUT_2_7,
  CRC_OUT_2_8,CRC_OUT_2_9,CRC_OUT_3_0,CRC_OUT_3_1,CRC_OUT_3_10,CRC_OUT_3_11,
  CRC_OUT_3_12,CRC_OUT_3_13,CRC_OUT_3_14,CRC_OUT_3_15,CRC_OUT_3_16,
  CRC_OUT_3_17,CRC_OUT_3_18,CRC_OUT_3_19,CRC_OUT_3_2,CRC_OUT_3_20,CRC_OUT_3_21,
  CRC_OUT_3_22,CRC_OUT_3_23,CRC_OUT_3_24,CRC_OUT_3_25,CRC_OUT_3_26,
  CRC_OUT_3_27,CRC_OUT_3_28,CRC_OUT_3_29,CRC_OUT_3_3,CRC_OUT_3_30,CRC_OUT_3_31,
  CRC_OUT_3_4,CRC_OUT_3_5,CRC_OUT_3_6,CRC_OUT_3_7,CRC_OUT_3_8,CRC_OUT_3_9,
  CRC_OUT_4_0,CRC_OUT_4_1,CRC_OUT_4_10,CRC_OUT_4_11,CRC_OUT_4_12,CRC_OUT_4_13,
  CRC_OUT_4_14,CRC_OUT_4_15,CRC_OUT_4_16,CRC_OUT_4_17,CRC_OUT_4_18,
  CRC_OUT_4_19,CRC_OUT_4_2,CRC_OUT_4_20,CRC_OUT_4_21,CRC_OUT_4_22,CRC_OUT_4_23,
  CRC_OUT_4_24,CRC_OUT_4_25,CRC_OUT_4_26,CRC_OUT_4_27,CRC_OUT_4_28,
  CRC_OUT_4_29,CRC_OUT_4_3,CRC_OUT_4_30,CRC_OUT_4_31,CRC_OUT_4_4,CRC_OUT_4_5,
  CRC_OUT_4_6,CRC_OUT_4_7,CRC_OUT_4_8,CRC_OUT_4_9,CRC_OUT_5_0,CRC_OUT_5_1,
  CRC_OUT_5_10,CRC_OUT_5_11,CRC_OUT_5_12,CRC_OUT_5_13,CRC_OUT_5_14,
  CRC_OUT_5_15,CRC_OUT_5_16,CRC_OUT_5_17,CRC_OUT_5_18,CRC_OUT_5_19,CRC_OUT_5_2,
  CRC_OUT_5_20,CRC_OUT_5_21,CRC_OUT_5_22,CRC_OUT_5_23,CRC_OUT_5_24,
  CRC_OUT_5_25,CRC_OUT_5_26,CRC_OUT_5_27,CRC_OUT_5_28,CRC_OUT_5_29,CRC_OUT_5_3,
  CRC_OUT_5_30,CRC_OUT_5_31,CRC_OUT_5_4,CRC_OUT_5_5,CRC_OUT_5_6,CRC_OUT_5_7,
  CRC_OUT_5_8,CRC_OUT_5_9,CRC_OUT_6_0,CRC_OUT_6_1,CRC_OUT_6_10,CRC_OUT_6_11,
  CRC_OUT_6_12,CRC_OUT_6_13,CRC_OUT_6_14,CRC_OUT_6_15,CRC_OUT_6_16,
  CRC_OUT_6_17,CRC_OUT_6_18,CRC_OUT_6_19,CRC_OUT_6_2,CRC_OUT_6_20,CRC_OUT_6_21,
  CRC_OUT_6_22,CRC_OUT_6_23,CRC_OUT_6_24,CRC_OUT_6_25,CRC_OUT_6_26,
  CRC_OUT_6_27,CRC_OUT_6_28,CRC_OUT_6_29,CRC_OUT_6_3,CRC_OUT_6_30,CRC_OUT_6_31,
  CRC_OUT_6_4,CRC_OUT_6_5,CRC_OUT_6_6,CRC_OUT_6_7,CRC_OUT_6_8,CRC_OUT_6_9,
  CRC_OUT_7_0,CRC_OUT_7_1,CRC_OUT_7_10,CRC_OUT_7_11,CRC_OUT_7_12,CRC_OUT_7_13,
  CRC_OUT_7_14,CRC_OUT_7_15,CRC_OUT_7_16,CRC_OUT_7_17,CRC_OUT_7_18,
  CRC_OUT_7_19,CRC_OUT_7_2,CRC_OUT_7_20,CRC_OUT_7_21,CRC_OUT_7_22,CRC_OUT_7_23,
  CRC_OUT_7_24,CRC_OUT_7_25,CRC_OUT_7_26,CRC_OUT_7_27,CRC_OUT_7_28,
  CRC_OUT_7_29,CRC_OUT_7_3,CRC_OUT_7_30,CRC_OUT_7_31,CRC_OUT_7_4,CRC_OUT_7_5,
  CRC_OUT_7_6,CRC_OUT_7_7,CRC_OUT_7_8,CRC_OUT_7_9,CRC_OUT_8_0,CRC_OUT_8_1,
  CRC_OUT_8_10,CRC_OUT_8_11,CRC_OUT_8_12,CRC_OUT_8_13,CRC_OUT_8_14,
  CRC_OUT_8_15,CRC_OUT_8_16,CRC_OUT_8_17,CRC_OUT_8_18,CRC_OUT_8_19,CRC_OUT_8_2,
  CRC_OUT_8_20,CRC_OUT_8_21,CRC_OUT_8_22,CRC_OUT_8_23,CRC_OUT_8_24,
  CRC_OUT_8_25,CRC_OUT_8_26,CRC_OUT_8_27,CRC_OUT_8_28,CRC_OUT_8_29,CRC_OUT_8_3,
  CRC_OUT_8_30,CRC_OUT_8_31,CRC_OUT_8_4,CRC_OUT_8_5,CRC_OUT_8_6,CRC_OUT_8_7,
  CRC_OUT_8_8,CRC_OUT_8_9,CRC_OUT_9_0,CRC_OUT_9_1,CRC_OUT_9_10,CRC_OUT_9_11,
  CRC_OUT_9_12,CRC_OUT_9_13,CRC_OUT_9_14,CRC_OUT_9_15,CRC_OUT_9_16,
  CRC_OUT_9_17,CRC_OUT_9_18,CRC_OUT_9_19,CRC_OUT_9_2,CRC_OUT_9_20,CRC_OUT_9_21,
  CRC_OUT_9_22,CRC_OUT_9_23,CRC_OUT_9_24,CRC_OUT_9_25,CRC_OUT_9_26,
  CRC_OUT_9_27,CRC_OUT_9_28,CRC_OUT_9_29,CRC_OUT_9_3,CRC_OUT_9_30,CRC_OUT_9_31,
  CRC_OUT_9_4,CRC_OUT_9_5,CRC_OUT_9_6,CRC_OUT_9_7,CRC_OUT_9_8,CRC_OUT_9_9,
  DATA_0_0,DATA_0_1,DATA_0_10,DATA_0_11,DATA_0_12,DATA_0_13,DATA_0_14,
  DATA_0_15,DATA_0_16,DATA_0_17,DATA_0_18,DATA_0_19,DATA_0_2,DATA_0_20,
  DATA_0_21,DATA_0_22,DATA_0_23,DATA_0_24,DATA_0_25,DATA_0_26,DATA_0_27,
  DATA_0_28,DATA_0_29,DATA_0_3,DATA_0_30,DATA_0_31,DATA_0_4,DATA_0_5,DATA_0_6,
  DATA_0_7,DATA_0_8,DATA_0_9,DATA_9_0,DATA_9_1,DATA_9_10,DATA_9_11,DATA_9_12,
  DATA_9_13,DATA_9_14,DATA_9_15,DATA_9_16,DATA_9_17,DATA_9_18,DATA_9_19,
  DATA_9_2,DATA_9_20,DATA_9_21,DATA_9_22,DATA_9_23,DATA_9_24,DATA_9_25,
  DATA_9_26,DATA_9_27,DATA_9_28,DATA_9_29,DATA_9_3,DATA_9_30,DATA_9_31,
  DATA_9_4,DATA_9_5,DATA_9_6,DATA_9_7,DATA_9_8,DATA_9_9,RESET,TM0,TM1);
input GND,VDD,CK,DATA_0_31,DATA_0_30,DATA_0_29,DATA_0_28,DATA_0_27,DATA_0_26,
  DATA_0_25,
  DATA_0_24,DATA_0_23,DATA_0_22,DATA_0_21,DATA_0_20,DATA_0_19,DATA_0_18,
  DATA_0_17,DATA_0_16,DATA_0_15,DATA_0_14,DATA_0_13,DATA_0_12,DATA_0_11,
  DATA_0_10,DATA_0_9,DATA_0_8,DATA_0_7,DATA_0_6,DATA_0_5,DATA_0_4,DATA_0_3,
  DATA_0_2,DATA_0_1,DATA_0_0,RESET,TM1,TM0;
output DATA_9_31,DATA_9_30,DATA_9_29,DATA_9_28,DATA_9_27,DATA_9_26,DATA_9_25,
  DATA_9_24,DATA_9_23,DATA_9_22,DATA_9_21,DATA_9_20,DATA_9_19,DATA_9_18,
  DATA_9_17,DATA_9_16,DATA_9_15,DATA_9_14,DATA_9_13,DATA_9_12,DATA_9_11,
  DATA_9_10,DATA_9_9,DATA_9_8,DATA_9_7,DATA_9_6,DATA_9_5,DATA_9_4,DATA_9_3,
  DATA_9_2,DATA_9_1,DATA_9_0,CRC_OUT_9_0,CRC_OUT_9_1,CRC_OUT_9_2,CRC_OUT_9_3,
  CRC_OUT_9_4,CRC_OUT_9_5,CRC_OUT_9_6,CRC_OUT_9_7,CRC_OUT_9_8,CRC_OUT_9_9,
  CRC_OUT_9_10,CRC_OUT_9_11,CRC_OUT_9_12,CRC_OUT_9_13,CRC_OUT_9_14,
  CRC_OUT_9_15,CRC_OUT_9_16,CRC_OUT_9_17,CRC_OUT_9_18,CRC_OUT_9_19,
  CRC_OUT_9_20,CRC_OUT_9_21,CRC_OUT_9_22,CRC_OUT_9_23,CRC_OUT_9_24,
  CRC_OUT_9_25,CRC_OUT_9_26,CRC_OUT_9_27,CRC_OUT_9_28,CRC_OUT_9_29,
  CRC_OUT_9_30,CRC_OUT_9_31,CRC_OUT_8_0,CRC_OUT_8_1,CRC_OUT_8_2,CRC_OUT_8_3,
  CRC_OUT_8_4,CRC_OUT_8_5,CRC_OUT_8_6,CRC_OUT_8_7,CRC_OUT_8_8,CRC_OUT_8_9,
  CRC_OUT_8_10,CRC_OUT_8_11,CRC_OUT_8_12,CRC_OUT_8_13,CRC_OUT_8_14,
  CRC_OUT_8_15,CRC_OUT_8_16,CRC_OUT_8_17,CRC_OUT_8_18,CRC_OUT_8_19,
  CRC_OUT_8_20,CRC_OUT_8_21,CRC_OUT_8_22,CRC_OUT_8_23,CRC_OUT_8_24,
  CRC_OUT_8_25,CRC_OUT_8_26,CRC_OUT_8_27,CRC_OUT_8_28,CRC_OUT_8_29,
  CRC_OUT_8_30,CRC_OUT_8_31,CRC_OUT_7_0,CRC_OUT_7_1,CRC_OUT_7_2,CRC_OUT_7_3,
  CRC_OUT_7_4,CRC_OUT_7_5,CRC_OUT_7_6,CRC_OUT_7_7,CRC_OUT_7_8,CRC_OUT_7_9,
  CRC_OUT_7_10,CRC_OUT_7_11,CRC_OUT_7_12,CRC_OUT_7_13,CRC_OUT_7_14,
  CRC_OUT_7_15,CRC_OUT_7_16,CRC_OUT_7_17,CRC_OUT_7_18,CRC_OUT_7_19,
  CRC_OUT_7_20,CRC_OUT_7_21,CRC_OUT_7_22,CRC_OUT_7_23,CRC_OUT_7_24,
  CRC_OUT_7_25,CRC_OUT_7_26,CRC_OUT_7_27,CRC_OUT_7_28,CRC_OUT_7_29,
  CRC_OUT_7_30,CRC_OUT_7_31,CRC_OUT_6_0,CRC_OUT_6_1,CRC_OUT_6_2,CRC_OUT_6_3,
  CRC_OUT_6_4,CRC_OUT_6_5,CRC_OUT_6_6,CRC_OUT_6_7,CRC_OUT_6_8,CRC_OUT_6_9,
  CRC_OUT_6_10,CRC_OUT_6_11,CRC_OUT_6_12,CRC_OUT_6_13,CRC_OUT_6_14,
  CRC_OUT_6_15,CRC_OUT_6_16,CRC_OUT_6_17,CRC_OUT_6_18,CRC_OUT_6_19,
  CRC_OUT_6_20,CRC_OUT_6_21,CRC_OUT_6_22,CRC_OUT_6_23,CRC_OUT_6_24,
  CRC_OUT_6_25,CRC_OUT_6_26,CRC_OUT_6_27,CRC_OUT_6_28,CRC_OUT_6_29,
  CRC_OUT_6_30,CRC_OUT_6_31,CRC_OUT_5_0,CRC_OUT_5_1,CRC_OUT_5_2,CRC_OUT_5_3,
  CRC_OUT_5_4,CRC_OUT_5_5,CRC_OUT_5_6,CRC_OUT_5_7,CRC_OUT_5_8,CRC_OUT_5_9,
  CRC_OUT_5_10,CRC_OUT_5_11,CRC_OUT_5_12,CRC_OUT_5_13,CRC_OUT_5_14,
  CRC_OUT_5_15,CRC_OUT_5_16,CRC_OUT_5_17,CRC_OUT_5_18,CRC_OUT_5_19,
  CRC_OUT_5_20,CRC_OUT_5_21,CRC_OUT_5_22,CRC_OUT_5_23,CRC_OUT_5_24,
  CRC_OUT_5_25,CRC_OUT_5_26,CRC_OUT_5_27,CRC_OUT_5_28,CRC_OUT_5_29,
  CRC_OUT_5_30,CRC_OUT_5_31,CRC_OUT_4_0,CRC_OUT_4_1,CRC_OUT_4_2,CRC_OUT_4_3,
  CRC_OUT_4_4,CRC_OUT_4_5,CRC_OUT_4_6,CRC_OUT_4_7,CRC_OUT_4_8,CRC_OUT_4_9,
  CRC_OUT_4_10,CRC_OUT_4_11,CRC_OUT_4_12,CRC_OUT_4_13,CRC_OUT_4_14,
  CRC_OUT_4_15,CRC_OUT_4_16,CRC_OUT_4_17,CRC_OUT_4_18,CRC_OUT_4_19,
  CRC_OUT_4_20,CRC_OUT_4_21,CRC_OUT_4_22,CRC_OUT_4_23,CRC_OUT_4_24,
  CRC_OUT_4_25,CRC_OUT_4_26,CRC_OUT_4_27,CRC_OUT_4_28,CRC_OUT_4_29,
  CRC_OUT_4_30,CRC_OUT_4_31,CRC_OUT_3_0,CRC_OUT_3_1,CRC_OUT_3_2,CRC_OUT_3_3,
  CRC_OUT_3_4,CRC_OUT_3_5,CRC_OUT_3_6,CRC_OUT_3_7,CRC_OUT_3_8,CRC_OUT_3_9,
  CRC_OUT_3_10,CRC_OUT_3_11,CRC_OUT_3_12,CRC_OUT_3_13,CRC_OUT_3_14,
  CRC_OUT_3_15,CRC_OUT_3_16,CRC_OUT_3_17,CRC_OUT_3_18,CRC_OUT_3_19,
  CRC_OUT_3_20,CRC_OUT_3_21,CRC_OUT_3_22,CRC_OUT_3_23,CRC_OUT_3_24,
  CRC_OUT_3_25,CRC_OUT_3_26,CRC_OUT_3_27,CRC_OUT_3_28,CRC_OUT_3_29,
  CRC_OUT_3_30,CRC_OUT_3_31,CRC_OUT_2_0,CRC_OUT_2_1,CRC_OUT_2_2,CRC_OUT_2_3,
  CRC_OUT_2_4,CRC_OUT_2_5,CRC_OUT_2_6,CRC_OUT_2_7,CRC_OUT_2_8,CRC_OUT_2_9,
  CRC_OUT_2_10,CRC_OUT_2_11,CRC_OUT_2_12,CRC_OUT_2_13,CRC_OUT_2_14,
  CRC_OUT_2_15,CRC_OUT_2_16,CRC_OUT_2_17,CRC_OUT_2_18,CRC_OUT_2_19,
  CRC_OUT_2_20,CRC_OUT_2_21,CRC_OUT_2_22,CRC_OUT_2_23,CRC_OUT_2_24,
  CRC_OUT_2_25,CRC_OUT_2_26,CRC_OUT_2_27,CRC_OUT_2_28,CRC_OUT_2_29,
  CRC_OUT_2_30,CRC_OUT_2_31,CRC_OUT_1_0,CRC_OUT_1_1,CRC_OUT_1_2,CRC_OUT_1_3,
  CRC_OUT_1_4,CRC_OUT_1_5,CRC_OUT_1_6,CRC_OUT_1_7,CRC_OUT_1_8,CRC_OUT_1_9,
  CRC_OUT_1_10,CRC_OUT_1_11,CRC_OUT_1_12,CRC_OUT_1_13,CRC_OUT_1_14,
  CRC_OUT_1_15,CRC_OUT_1_16,CRC_OUT_1_17,CRC_OUT_1_18,CRC_OUT_1_19,
  CRC_OUT_1_20,CRC_OUT_1_21,CRC_OUT_1_22,CRC_OUT_1_23,CRC_OUT_1_24,
  CRC_OUT_1_25,CRC_OUT_1_26,CRC_OUT_1_27,CRC_OUT_1_28,CRC_OUT_1_29,
  CRC_OUT_1_30,CRC_OUT_1_31;

  wire WX485,WX484,WX487,WX486,WX489,WX488,WX491,WX490,WX493,WX492,WX495,WX494,
    WX497,WX496,WX499,WX498,WX501,WX500,WX503,WX502,WX505,WX504,WX507,WX506,
    WX509,WX508,WX511,WX510,WX513,WX512,WX515,WX514,WX517,WX516,WX519,WX518,
    WX521,WX520,WX523,WX522,WX525,WX524,WX527,WX526,WX529,WX528,WX531,WX530,
    WX533,WX532,WX535,WX534,WX537,WX536,WX539,WX538,WX541,WX540,WX543,WX542,
    WX545,WX544,WX547,WX546,WX645,WX644,WX647,WX646,WX649,WX648,WX651,WX650,
    WX653,WX652,WX655,WX654,WX657,WX656,WX659,WX658,WX661,WX660,WX663,WX662,
    WX665,WX664,WX667,WX666,WX669,WX668,WX671,WX670,WX673,WX672,WX675,WX674,
    WX677,WX676,WX679,WX678,WX681,WX680,WX683,WX682,WX685,WX684,WX687,WX686,
    WX689,WX688,WX691,WX690,WX693,WX692,WX695,WX694,WX697,WX696,WX699,WX698,
    WX701,WX700,WX703,WX702,WX705,WX704,WX707,WX706,WX709,WX708,WX711,WX710,
    WX713,WX712,WX715,WX714,WX717,WX716,WX719,WX718,WX721,WX720,WX723,WX722,
    WX725,WX724,WX727,WX726,WX729,WX728,WX731,WX730,WX733,WX732,WX735,WX734,
    WX737,WX736,WX739,WX738,WX741,WX740,WX743,WX742,WX745,WX744,WX747,WX746,
    WX749,WX748,WX751,WX750,WX753,WX752,WX755,WX754,WX757,WX756,WX759,WX758,
    WX761,WX760,WX763,WX762,WX765,WX764,WX767,WX766,WX769,WX768,WX771,WX770,
    WX773,WX772,WX775,WX774,WX777,WX776,WX779,WX778,WX781,WX780,WX783,WX782,
    WX785,WX784,WX787,WX786,WX789,WX788,WX791,WX790,WX793,WX792,WX795,WX794,
    WX797,WX796,WX799,WX798,WX801,WX800,WX803,WX802,WX805,WX804,WX807,WX806,
    WX809,WX808,WX811,WX810,WX813,WX812,WX815,WX814,WX817,WX816,WX819,WX818,
    WX821,WX820,WX823,WX822,WX825,WX824,WX827,WX826,WX829,WX828,WX831,WX830,
    WX833,WX832,WX835,WX834,WX837,WX836,WX839,WX838,WX841,WX840,WX843,WX842,
    WX845,WX844,WX847,WX846,WX849,WX848,WX851,WX850,WX853,WX852,WX855,WX854,
    WX857,WX856,WX859,WX858,WX861,WX860,WX863,WX862,WX865,WX864,WX867,WX866,
    WX869,WX868,WX871,WX870,WX873,WX872,WX875,WX874,WX877,WX876,WX879,WX878,
    WX881,WX880,WX883,WX882,WX885,WX884,WX887,WX886,WX889,WX888,WX891,WX890,
    WX893,WX892,WX895,WX894,WX897,WX896,WX899,WX898,WX1264,WX1266,WX1268,
    WX1270,WX1272,WX1274,WX1276,WX1278,WX1280,WX1282,WX1284,WX1286,WX1288,
    WX1290,WX1292,WX1294,WX1296,WX1298,WX1300,WX1302,WX1304,WX1306,WX1308,
    WX1310,WX1312,WX1314,WX1316,WX1318,WX1320,WX1322,WX1324,WX1326,WX1778,
    WX1777,WX1780,WX1779,WX1782,WX1781,WX1784,WX1783,WX1786,WX1785,WX1788,
    WX1787,WX1790,WX1789,WX1792,WX1791,WX1794,WX1793,WX1796,WX1795,WX1798,
    WX1797,WX1800,WX1799,WX1802,WX1801,WX1804,WX1803,WX1806,WX1805,WX1808,
    WX1807,WX1810,WX1809,WX1812,WX1811,WX1814,WX1813,WX1816,WX1815,WX1818,
    WX1817,WX1820,WX1819,WX1822,WX1821,WX1824,WX1823,WX1826,WX1825,WX1828,
    WX1827,WX1830,WX1829,WX1832,WX1831,WX1834,WX1833,WX1836,WX1835,WX1838,
    WX1837,WX1840,WX1839,WX1938,WX1937,WX1940,WX1939,WX1942,WX1941,WX1944,
    WX1943,WX1946,WX1945,WX1948,WX1947,WX1950,WX1949,WX1952,WX1951,WX1954,
    WX1953,WX1956,WX1955,WX1958,WX1957,WX1960,WX1959,WX1962,WX1961,WX1964,
    WX1963,WX1966,WX1965,WX1968,WX1967,WX1970,WX1969,WX1972,WX1971,WX1974,
    WX1973,WX1976,WX1975,WX1978,WX1977,WX1980,WX1979,WX1982,WX1981,WX1984,
    WX1983,WX1986,WX1985,WX1988,WX1987,WX1990,WX1989,WX1992,WX1991,WX1994,
    WX1993,WX1996,WX1995,WX1998,WX1997,WX2000,WX1999,WX2002,WX2001,WX2004,
    WX2003,WX2006,WX2005,WX2008,WX2007,WX2010,WX2009,WX2012,WX2011,WX2014,
    WX2013,WX2016,WX2015,WX2018,WX2017,WX2020,WX2019,WX2022,WX2021,WX2024,
    WX2023,WX2026,WX2025,WX2028,WX2027,WX2030,WX2029,WX2032,WX2031,WX2034,
    WX2033,WX2036,WX2035,WX2038,WX2037,WX2040,WX2039,WX2042,WX2041,WX2044,
    WX2043,WX2046,WX2045,WX2048,WX2047,WX2050,WX2049,WX2052,WX2051,WX2054,
    WX2053,WX2056,WX2055,WX2058,WX2057,WX2060,WX2059,WX2062,WX2061,WX2064,
    WX2063,WX2066,WX2065,WX2068,WX2067,WX2070,WX2069,WX2072,WX2071,WX2074,
    WX2073,WX2076,WX2075,WX2078,WX2077,WX2080,WX2079,WX2082,WX2081,WX2084,
    WX2083,WX2086,WX2085,WX2088,WX2087,WX2090,WX2089,WX2092,WX2091,WX2094,
    WX2093,WX2096,WX2095,WX2098,WX2097,WX2100,WX2099,WX2102,WX2101,WX2104,
    WX2103,WX2106,WX2105,WX2108,WX2107,WX2110,WX2109,WX2112,WX2111,WX2114,
    WX2113,WX2116,WX2115,WX2118,WX2117,WX2120,WX2119,WX2122,WX2121,WX2124,
    WX2123,WX2126,WX2125,WX2128,WX2127,WX2130,WX2129,WX2132,WX2131,WX2134,
    WX2133,WX2136,WX2135,WX2138,WX2137,WX2140,WX2139,WX2142,WX2141,WX2144,
    WX2143,WX2146,WX2145,WX2148,WX2147,WX2150,WX2149,WX2152,WX2151,WX2154,
    WX2153,WX2156,WX2155,WX2158,WX2157,WX2160,WX2159,WX2162,WX2161,WX2164,
    WX2163,WX2166,WX2165,WX2168,WX2167,WX2170,WX2169,WX2172,WX2171,WX2174,
    WX2173,WX2176,WX2175,WX2178,WX2177,WX2180,WX2179,WX2182,WX2181,WX2184,
    WX2183,WX2186,WX2185,WX2188,WX2187,WX2190,WX2189,WX2192,WX2191,WX2557,
    WX2559,WX2561,WX2563,WX2565,WX2567,WX2569,WX2571,WX2573,WX2575,WX2577,
    WX2579,WX2581,WX2583,WX2585,WX2587,WX2589,WX2591,WX2593,WX2595,WX2597,
    WX2599,WX2601,WX2603,WX2605,WX2607,WX2609,WX2611,WX2613,WX2615,WX2617,
    WX2619,WX3071,WX3070,WX3073,WX3072,WX3075,WX3074,WX3077,WX3076,WX3079,
    WX3078,WX3081,WX3080,WX3083,WX3082,WX3085,WX3084,WX3087,WX3086,WX3089,
    WX3088,WX3091,WX3090,WX3093,WX3092,WX3095,WX3094,WX3097,WX3096,WX3099,
    WX3098,WX3101,WX3100,WX3103,WX3102,WX3105,WX3104,WX3107,WX3106,WX3109,
    WX3108,WX3111,WX3110,WX3113,WX3112,WX3115,WX3114,WX3117,WX3116,WX3119,
    WX3118,WX3121,WX3120,WX3123,WX3122,WX3125,WX3124,WX3127,WX3126,WX3129,
    WX3128,WX3131,WX3130,WX3133,WX3132,WX3231,WX3230,WX3233,WX3232,WX3235,
    WX3234,WX3237,WX3236,WX3239,WX3238,WX3241,WX3240,WX3243,WX3242,WX3245,
    WX3244,WX3247,WX3246,WX3249,WX3248,WX3251,WX3250,WX3253,WX3252,WX3255,
    WX3254,WX3257,WX3256,WX3259,WX3258,WX3261,WX3260,WX3263,WX3262,WX3265,
    WX3264,WX3267,WX3266,WX3269,WX3268,WX3271,WX3270,WX3273,WX3272,WX3275,
    WX3274,WX3277,WX3276,WX3279,WX3278,WX3281,WX3280,WX3283,WX3282,WX3285,
    WX3284,WX3287,WX3286,WX3289,WX3288,WX3291,WX3290,WX3293,WX3292,WX3295,
    WX3294,WX3297,WX3296,WX3299,WX3298,WX3301,WX3300,WX3303,WX3302,WX3305,
    WX3304,WX3307,WX3306,WX3309,WX3308,WX3311,WX3310,WX3313,WX3312,WX3315,
    WX3314,WX3317,WX3316,WX3319,WX3318,WX3321,WX3320,WX3323,WX3322,WX3325,
    WX3324,WX3327,WX3326,WX3329,WX3328,WX3331,WX3330,WX3333,WX3332,WX3335,
    WX3334,WX3337,WX3336,WX3339,WX3338,WX3341,WX3340,WX3343,WX3342,WX3345,
    WX3344,WX3347,WX3346,WX3349,WX3348,WX3351,WX3350,WX3353,WX3352,WX3355,
    WX3354,WX3357,WX3356,WX3359,WX3358,WX3361,WX3360,WX3363,WX3362,WX3365,
    WX3364,WX3367,WX3366,WX3369,WX3368,WX3371,WX3370,WX3373,WX3372,WX3375,
    WX3374,WX3377,WX3376,WX3379,WX3378,WX3381,WX3380,WX3383,WX3382,WX3385,
    WX3384,WX3387,WX3386,WX3389,WX3388,WX3391,WX3390,WX3393,WX3392,WX3395,
    WX3394,WX3397,WX3396,WX3399,WX3398,WX3401,WX3400,WX3403,WX3402,WX3405,
    WX3404,WX3407,WX3406,WX3409,WX3408,WX3411,WX3410,WX3413,WX3412,WX3415,
    WX3414,WX3417,WX3416,WX3419,WX3418,WX3421,WX3420,WX3423,WX3422,WX3425,
    WX3424,WX3427,WX3426,WX3429,WX3428,WX3431,WX3430,WX3433,WX3432,WX3435,
    WX3434,WX3437,WX3436,WX3439,WX3438,WX3441,WX3440,WX3443,WX3442,WX3445,
    WX3444,WX3447,WX3446,WX3449,WX3448,WX3451,WX3450,WX3453,WX3452,WX3455,
    WX3454,WX3457,WX3456,WX3459,WX3458,WX3461,WX3460,WX3463,WX3462,WX3465,
    WX3464,WX3467,WX3466,WX3469,WX3468,WX3471,WX3470,WX3473,WX3472,WX3475,
    WX3474,WX3477,WX3476,WX3479,WX3478,WX3481,WX3480,WX3483,WX3482,WX3485,
    WX3484,WX3850,WX3852,WX3854,WX3856,WX3858,WX3860,WX3862,WX3864,WX3866,
    WX3868,WX3870,WX3872,WX3874,WX3876,WX3878,WX3880,WX3882,WX3884,WX3886,
    WX3888,WX3890,WX3892,WX3894,WX3896,WX3898,WX3900,WX3902,WX3904,WX3906,
    WX3908,WX3910,WX3912,WX4364,WX4363,WX4366,WX4365,WX4368,WX4367,WX4370,
    WX4369,WX4372,WX4371,WX4374,WX4373,WX4376,WX4375,WX4378,WX4377,WX4380,
    WX4379,WX4382,WX4381,WX4384,WX4383,WX4386,WX4385,WX4388,WX4387,WX4390,
    WX4389,WX4392,WX4391,WX4394,WX4393,WX4396,WX4395,WX4398,WX4397,WX4400,
    WX4399,WX4402,WX4401,WX4404,WX4403,WX4406,WX4405,WX4408,WX4407,WX4410,
    WX4409,WX4412,WX4411,WX4414,WX4413,WX4416,WX4415,WX4418,WX4417,WX4420,
    WX4419,WX4422,WX4421,WX4424,WX4423,WX4426,WX4425,WX4524,WX4523,WX4526,
    WX4525,WX4528,WX4527,WX4530,WX4529,WX4532,WX4531,WX4534,WX4533,WX4536,
    WX4535,WX4538,WX4537,WX4540,WX4539,WX4542,WX4541,WX4544,WX4543,WX4546,
    WX4545,WX4548,WX4547,WX4550,WX4549,WX4552,WX4551,WX4554,WX4553,WX4556,
    WX4555,WX4558,WX4557,WX4560,WX4559,WX4562,WX4561,WX4564,WX4563,WX4566,
    WX4565,WX4568,WX4567,WX4570,WX4569,WX4572,WX4571,WX4574,WX4573,WX4576,
    WX4575,WX4578,WX4577,WX4580,WX4579,WX4582,WX4581,WX4584,WX4583,WX4586,
    WX4585,WX4588,WX4587,WX4590,WX4589,WX4592,WX4591,WX4594,WX4593,WX4596,
    WX4595,WX4598,WX4597,WX4600,WX4599,WX4602,WX4601,WX4604,WX4603,WX4606,
    WX4605,WX4608,WX4607,WX4610,WX4609,WX4612,WX4611,WX4614,WX4613,WX4616,
    WX4615,WX4618,WX4617,WX4620,WX4619,WX4622,WX4621,WX4624,WX4623,WX4626,
    WX4625,WX4628,WX4627,WX4630,WX4629,WX4632,WX4631,WX4634,WX4633,WX4636,
    WX4635,WX4638,WX4637,WX4640,WX4639,WX4642,WX4641,WX4644,WX4643,WX4646,
    WX4645,WX4648,WX4647,WX4650,WX4649,WX4652,WX4651,WX4654,WX4653,WX4656,
    WX4655,WX4658,WX4657,WX4660,WX4659,WX4662,WX4661,WX4664,WX4663,WX4666,
    WX4665,WX4668,WX4667,WX4670,WX4669,WX4672,WX4671,WX4674,WX4673,WX4676,
    WX4675,WX4678,WX4677,WX4680,WX4679,WX4682,WX4681,WX4684,WX4683,WX4686,
    WX4685,WX4688,WX4687,WX4690,WX4689,WX4692,WX4691,WX4694,WX4693,WX4696,
    WX4695,WX4698,WX4697,WX4700,WX4699,WX4702,WX4701,WX4704,WX4703,WX4706,
    WX4705,WX4708,WX4707,WX4710,WX4709,WX4712,WX4711,WX4714,WX4713,WX4716,
    WX4715,WX4718,WX4717,WX4720,WX4719,WX4722,WX4721,WX4724,WX4723,WX4726,
    WX4725,WX4728,WX4727,WX4730,WX4729,WX4732,WX4731,WX4734,WX4733,WX4736,
    WX4735,WX4738,WX4737,WX4740,WX4739,WX4742,WX4741,WX4744,WX4743,WX4746,
    WX4745,WX4748,WX4747,WX4750,WX4749,WX4752,WX4751,WX4754,WX4753,WX4756,
    WX4755,WX4758,WX4757,WX4760,WX4759,WX4762,WX4761,WX4764,WX4763,WX4766,
    WX4765,WX4768,WX4767,WX4770,WX4769,WX4772,WX4771,WX4774,WX4773,WX4776,
    WX4775,WX4778,WX4777,WX5143,WX5145,WX5147,WX5149,WX5151,WX5153,WX5155,
    WX5157,WX5159,WX5161,WX5163,WX5165,WX5167,WX5169,WX5171,WX5173,WX5175,
    WX5177,WX5179,WX5181,WX5183,WX5185,WX5187,WX5189,WX5191,WX5193,WX5195,
    WX5197,WX5199,WX5201,WX5203,WX5205,WX5657,WX5656,WX5659,WX5658,WX5661,
    WX5660,WX5663,WX5662,WX5665,WX5664,WX5667,WX5666,WX5669,WX5668,WX5671,
    WX5670,WX5673,WX5672,WX5675,WX5674,WX5677,WX5676,WX5679,WX5678,WX5681,
    WX5680,WX5683,WX5682,WX5685,WX5684,WX5687,WX5686,WX5689,WX5688,WX5691,
    WX5690,WX5693,WX5692,WX5695,WX5694,WX5697,WX5696,WX5699,WX5698,WX5701,
    WX5700,WX5703,WX5702,WX5705,WX5704,WX5707,WX5706,WX5709,WX5708,WX5711,
    WX5710,WX5713,WX5712,WX5715,WX5714,WX5717,WX5716,WX5719,WX5718,WX5817,
    WX5816,WX5819,WX5818,WX5821,WX5820,WX5823,WX5822,WX5825,WX5824,WX5827,
    WX5826,WX5829,WX5828,WX5831,WX5830,WX5833,WX5832,WX5835,WX5834,WX5837,
    WX5836,WX5839,WX5838,WX5841,WX5840,WX5843,WX5842,WX5845,WX5844,WX5847,
    WX5846,WX5849,WX5848,WX5851,WX5850,WX5853,WX5852,WX5855,WX5854,WX5857,
    WX5856,WX5859,WX5858,WX5861,WX5860,WX5863,WX5862,WX5865,WX5864,WX5867,
    WX5866,WX5869,WX5868,WX5871,WX5870,WX5873,WX5872,WX5875,WX5874,WX5877,
    WX5876,WX5879,WX5878,WX5881,WX5880,WX5883,WX5882,WX5885,WX5884,WX5887,
    WX5886,WX5889,WX5888,WX5891,WX5890,WX5893,WX5892,WX5895,WX5894,WX5897,
    WX5896,WX5899,WX5898,WX5901,WX5900,WX5903,WX5902,WX5905,WX5904,WX5907,
    WX5906,WX5909,WX5908,WX5911,WX5910,WX5913,WX5912,WX5915,WX5914,WX5917,
    WX5916,WX5919,WX5918,WX5921,WX5920,WX5923,WX5922,WX5925,WX5924,WX5927,
    WX5926,WX5929,WX5928,WX5931,WX5930,WX5933,WX5932,WX5935,WX5934,WX5937,
    WX5936,WX5939,WX5938,WX5941,WX5940,WX5943,WX5942,WX5945,WX5944,WX5947,
    WX5946,WX5949,WX5948,WX5951,WX5950,WX5953,WX5952,WX5955,WX5954,WX5957,
    WX5956,WX5959,WX5958,WX5961,WX5960,WX5963,WX5962,WX5965,WX5964,WX5967,
    WX5966,WX5969,WX5968,WX5971,WX5970,WX5973,WX5972,WX5975,WX5974,WX5977,
    WX5976,WX5979,WX5978,WX5981,WX5980,WX5983,WX5982,WX5985,WX5984,WX5987,
    WX5986,WX5989,WX5988,WX5991,WX5990,WX5993,WX5992,WX5995,WX5994,WX5997,
    WX5996,WX5999,WX5998,WX6001,WX6000,WX6003,WX6002,WX6005,WX6004,WX6007,
    WX6006,WX6009,WX6008,WX6011,WX6010,WX6013,WX6012,WX6015,WX6014,WX6017,
    WX6016,WX6019,WX6018,WX6021,WX6020,WX6023,WX6022,WX6025,WX6024,WX6027,
    WX6026,WX6029,WX6028,WX6031,WX6030,WX6033,WX6032,WX6035,WX6034,WX6037,
    WX6036,WX6039,WX6038,WX6041,WX6040,WX6043,WX6042,WX6045,WX6044,WX6047,
    WX6046,WX6049,WX6048,WX6051,WX6050,WX6053,WX6052,WX6055,WX6054,WX6057,
    WX6056,WX6059,WX6058,WX6061,WX6060,WX6063,WX6062,WX6065,WX6064,WX6067,
    WX6066,WX6069,WX6068,WX6071,WX6070,WX6436,WX6438,WX6440,WX6442,WX6444,
    WX6446,WX6448,WX6450,WX6452,WX6454,WX6456,WX6458,WX6460,WX6462,WX6464,
    WX6466,WX6468,WX6470,WX6472,WX6474,WX6476,WX6478,WX6480,WX6482,WX6484,
    WX6486,WX6488,WX6490,WX6492,WX6494,WX6496,WX6498,WX6950,WX6949,WX6952,
    WX6951,WX6954,WX6953,WX6956,WX6955,WX6958,WX6957,WX6960,WX6959,WX6962,
    WX6961,WX6964,WX6963,WX6966,WX6965,WX6968,WX6967,WX6970,WX6969,WX6972,
    WX6971,WX6974,WX6973,WX6976,WX6975,WX6978,WX6977,WX6980,WX6979,WX6982,
    WX6981,WX6984,WX6983,WX6986,WX6985,WX6988,WX6987,WX6990,WX6989,WX6992,
    WX6991,WX6994,WX6993,WX6996,WX6995,WX6998,WX6997,WX7000,WX6999,WX7002,
    WX7001,WX7004,WX7003,WX7006,WX7005,WX7008,WX7007,WX7010,WX7009,WX7012,
    WX7011,WX7110,WX7109,WX7112,WX7111,WX7114,WX7113,WX7116,WX7115,WX7118,
    WX7117,WX7120,WX7119,WX7122,WX7121,WX7124,WX7123,WX7126,WX7125,WX7128,
    WX7127,WX7130,WX7129,WX7132,WX7131,WX7134,WX7133,WX7136,WX7135,WX7138,
    WX7137,WX7140,WX7139,WX7142,WX7141,WX7144,WX7143,WX7146,WX7145,WX7148,
    WX7147,WX7150,WX7149,WX7152,WX7151,WX7154,WX7153,WX7156,WX7155,WX7158,
    WX7157,WX7160,WX7159,WX7162,WX7161,WX7164,WX7163,WX7166,WX7165,WX7168,
    WX7167,WX7170,WX7169,WX7172,WX7171,WX7174,WX7173,WX7176,WX7175,WX7178,
    WX7177,WX7180,WX7179,WX7182,WX7181,WX7184,WX7183,WX7186,WX7185,WX7188,
    WX7187,WX7190,WX7189,WX7192,WX7191,WX7194,WX7193,WX7196,WX7195,WX7198,
    WX7197,WX7200,WX7199,WX7202,WX7201,WX7204,WX7203,WX7206,WX7205,WX7208,
    WX7207,WX7210,WX7209,WX7212,WX7211,WX7214,WX7213,WX7216,WX7215,WX7218,
    WX7217,WX7220,WX7219,WX7222,WX7221,WX7224,WX7223,WX7226,WX7225,WX7228,
    WX7227,WX7230,WX7229,WX7232,WX7231,WX7234,WX7233,WX7236,WX7235,WX7238,
    WX7237,WX7240,WX7239,WX7242,WX7241,WX7244,WX7243,WX7246,WX7245,WX7248,
    WX7247,WX7250,WX7249,WX7252,WX7251,WX7254,WX7253,WX7256,WX7255,WX7258,
    WX7257,WX7260,WX7259,WX7262,WX7261,WX7264,WX7263,WX7266,WX7265,WX7268,
    WX7267,WX7270,WX7269,WX7272,WX7271,WX7274,WX7273,WX7276,WX7275,WX7278,
    WX7277,WX7280,WX7279,WX7282,WX7281,WX7284,WX7283,WX7286,WX7285,WX7288,
    WX7287,WX7290,WX7289,WX7292,WX7291,WX7294,WX7293,WX7296,WX7295,WX7298,
    WX7297,WX7300,WX7299,WX7302,WX7301,WX7304,WX7303,WX7306,WX7305,WX7308,
    WX7307,WX7310,WX7309,WX7312,WX7311,WX7314,WX7313,WX7316,WX7315,WX7318,
    WX7317,WX7320,WX7319,WX7322,WX7321,WX7324,WX7323,WX7326,WX7325,WX7328,
    WX7327,WX7330,WX7329,WX7332,WX7331,WX7334,WX7333,WX7336,WX7335,WX7338,
    WX7337,WX7340,WX7339,WX7342,WX7341,WX7344,WX7343,WX7346,WX7345,WX7348,
    WX7347,WX7350,WX7349,WX7352,WX7351,WX7354,WX7353,WX7356,WX7355,WX7358,
    WX7357,WX7360,WX7359,WX7362,WX7361,WX7364,WX7363,WX7729,WX7731,WX7733,
    WX7735,WX7737,WX7739,WX7741,WX7743,WX7745,WX7747,WX7749,WX7751,WX7753,
    WX7755,WX7757,WX7759,WX7761,WX7763,WX7765,WX7767,WX7769,WX7771,WX7773,
    WX7775,WX7777,WX7779,WX7781,WX7783,WX7785,WX7787,WX7789,WX7791,WX8243,
    WX8242,WX8245,WX8244,WX8247,WX8246,WX8249,WX8248,WX8251,WX8250,WX8253,
    WX8252,WX8255,WX8254,WX8257,WX8256,WX8259,WX8258,WX8261,WX8260,WX8263,
    WX8262,WX8265,WX8264,WX8267,WX8266,WX8269,WX8268,WX8271,WX8270,WX8273,
    WX8272,WX8275,WX8274,WX8277,WX8276,WX8279,WX8278,WX8281,WX8280,WX8283,
    WX8282,WX8285,WX8284,WX8287,WX8286,WX8289,WX8288,WX8291,WX8290,WX8293,
    WX8292,WX8295,WX8294,WX8297,WX8296,WX8299,WX8298,WX8301,WX8300,WX8303,
    WX8302,WX8305,WX8304,WX8403,WX8402,WX8405,WX8404,WX8407,WX8406,WX8409,
    WX8408,WX8411,WX8410,WX8413,WX8412,WX8415,WX8414,WX8417,WX8416,WX8419,
    WX8418,WX8421,WX8420,WX8423,WX8422,WX8425,WX8424,WX8427,WX8426,WX8429,
    WX8428,WX8431,WX8430,WX8433,WX8432,WX8435,WX8434,WX8437,WX8436,WX8439,
    WX8438,WX8441,WX8440,WX8443,WX8442,WX8445,WX8444,WX8447,WX8446,WX8449,
    WX8448,WX8451,WX8450,WX8453,WX8452,WX8455,WX8454,WX8457,WX8456,WX8459,
    WX8458,WX8461,WX8460,WX8463,WX8462,WX8465,WX8464,WX8467,WX8466,WX8469,
    WX8468,WX8471,WX8470,WX8473,WX8472,WX8475,WX8474,WX8477,WX8476,WX8479,
    WX8478,WX8481,WX8480,WX8483,WX8482,WX8485,WX8484,WX8487,WX8486,WX8489,
    WX8488,WX8491,WX8490,WX8493,WX8492,WX8495,WX8494,WX8497,WX8496,WX8499,
    WX8498,WX8501,WX8500,WX8503,WX8502,WX8505,WX8504,WX8507,WX8506,WX8509,
    WX8508,WX8511,WX8510,WX8513,WX8512,WX8515,WX8514,WX8517,WX8516,WX8519,
    WX8518,WX8521,WX8520,WX8523,WX8522,WX8525,WX8524,WX8527,WX8526,WX8529,
    WX8528,WX8531,WX8530,WX8533,WX8532,WX8535,WX8534,WX8537,WX8536,WX8539,
    WX8538,WX8541,WX8540,WX8543,WX8542,WX8545,WX8544,WX8547,WX8546,WX8549,
    WX8548,WX8551,WX8550,WX8553,WX8552,WX8555,WX8554,WX8557,WX8556,WX8559,
    WX8558,WX8561,WX8560,WX8563,WX8562,WX8565,WX8564,WX8567,WX8566,WX8569,
    WX8568,WX8571,WX8570,WX8573,WX8572,WX8575,WX8574,WX8577,WX8576,WX8579,
    WX8578,WX8581,WX8580,WX8583,WX8582,WX8585,WX8584,WX8587,WX8586,WX8589,
    WX8588,WX8591,WX8590,WX8593,WX8592,WX8595,WX8594,WX8597,WX8596,WX8599,
    WX8598,WX8601,WX8600,WX8603,WX8602,WX8605,WX8604,WX8607,WX8606,WX8609,
    WX8608,WX8611,WX8610,WX8613,WX8612,WX8615,WX8614,WX8617,WX8616,WX8619,
    WX8618,WX8621,WX8620,WX8623,WX8622,WX8625,WX8624,WX8627,WX8626,WX8629,
    WX8628,WX8631,WX8630,WX8633,WX8632,WX8635,WX8634,WX8637,WX8636,WX8639,
    WX8638,WX8641,WX8640,WX8643,WX8642,WX8645,WX8644,WX8647,WX8646,WX8649,
    WX8648,WX8651,WX8650,WX8653,WX8652,WX8655,WX8654,WX8657,WX8656,WX9022,
    WX9024,WX9026,WX9028,WX9030,WX9032,WX9034,WX9036,WX9038,WX9040,WX9042,
    WX9044,WX9046,WX9048,WX9050,WX9052,WX9054,WX9056,WX9058,WX9060,WX9062,
    WX9064,WX9066,WX9068,WX9070,WX9072,WX9074,WX9076,WX9078,WX9080,WX9082,
    WX9084,WX9536,WX9535,WX9538,WX9537,WX9540,WX9539,WX9542,WX9541,WX9544,
    WX9543,WX9546,WX9545,WX9548,WX9547,WX9550,WX9549,WX9552,WX9551,WX9554,
    WX9553,WX9556,WX9555,WX9558,WX9557,WX9560,WX9559,WX9562,WX9561,WX9564,
    WX9563,WX9566,WX9565,WX9568,WX9567,WX9570,WX9569,WX9572,WX9571,WX9574,
    WX9573,WX9576,WX9575,WX9578,WX9577,WX9580,WX9579,WX9582,WX9581,WX9584,
    WX9583,WX9586,WX9585,WX9588,WX9587,WX9590,WX9589,WX9592,WX9591,WX9594,
    WX9593,WX9596,WX9595,WX9598,WX9597,WX9696,WX9695,WX9698,WX9697,WX9700,
    WX9699,WX9702,WX9701,WX9704,WX9703,WX9706,WX9705,WX9708,WX9707,WX9710,
    WX9709,WX9712,WX9711,WX9714,WX9713,WX9716,WX9715,WX9718,WX9717,WX9720,
    WX9719,WX9722,WX9721,WX9724,WX9723,WX9726,WX9725,WX9728,WX9727,WX9730,
    WX9729,WX9732,WX9731,WX9734,WX9733,WX9736,WX9735,WX9738,WX9737,WX9740,
    WX9739,WX9742,WX9741,WX9744,WX9743,WX9746,WX9745,WX9748,WX9747,WX9750,
    WX9749,WX9752,WX9751,WX9754,WX9753,WX9756,WX9755,WX9758,WX9757,WX9760,
    WX9759,WX9762,WX9761,WX9764,WX9763,WX9766,WX9765,WX9768,WX9767,WX9770,
    WX9769,WX9772,WX9771,WX9774,WX9773,WX9776,WX9775,WX9778,WX9777,WX9780,
    WX9779,WX9782,WX9781,WX9784,WX9783,WX9786,WX9785,WX9788,WX9787,WX9790,
    WX9789,WX9792,WX9791,WX9794,WX9793,WX9796,WX9795,WX9798,WX9797,WX9800,
    WX9799,WX9802,WX9801,WX9804,WX9803,WX9806,WX9805,WX9808,WX9807,WX9810,
    WX9809,WX9812,WX9811,WX9814,WX9813,WX9816,WX9815,WX9818,WX9817,WX9820,
    WX9819,WX9822,WX9821,WX9824,WX9823,WX9826,WX9825,WX9828,WX9827,WX9830,
    WX9829,WX9832,WX9831,WX9834,WX9833,WX9836,WX9835,WX9838,WX9837,WX9840,
    WX9839,WX9842,WX9841,WX9844,WX9843,WX9846,WX9845,WX9848,WX9847,WX9850,
    WX9849,WX9852,WX9851,WX9854,WX9853,WX9856,WX9855,WX9858,WX9857,WX9860,
    WX9859,WX9862,WX9861,WX9864,WX9863,WX9866,WX9865,WX9868,WX9867,WX9870,
    WX9869,WX9872,WX9871,WX9874,WX9873,WX9876,WX9875,WX9878,WX9877,WX9880,
    WX9879,WX9882,WX9881,WX9884,WX9883,WX9886,WX9885,WX9888,WX9887,WX9890,
    WX9889,WX9892,WX9891,WX9894,WX9893,WX9896,WX9895,WX9898,WX9897,WX9900,
    WX9899,WX9902,WX9901,WX9904,WX9903,WX9906,WX9905,WX9908,WX9907,WX9910,
    WX9909,WX9912,WX9911,WX9914,WX9913,WX9916,WX9915,WX9918,WX9917,WX9920,
    WX9919,WX9922,WX9921,WX9924,WX9923,WX9926,WX9925,WX9928,WX9927,WX9930,
    WX9929,WX9932,WX9931,WX9934,WX9933,WX9936,WX9935,WX9938,WX9937,WX9940,
    WX9939,WX9942,WX9941,WX9944,WX9943,WX9946,WX9945,WX9948,WX9947,WX9950,
    WX9949,WX10315,WX10317,WX10319,WX10321,WX10323,WX10325,WX10327,WX10329,
    WX10331,WX10333,WX10335,WX10337,WX10339,WX10341,WX10343,WX10345,WX10347,
    WX10349,WX10351,WX10353,WX10355,WX10357,WX10359,WX10361,WX10363,WX10365,
    WX10367,WX10369,WX10371,WX10373,WX10375,WX10377,WX10829,WX10828,WX10831,
    WX10830,WX10833,WX10832,WX10835,WX10834,WX10837,WX10836,WX10839,WX10838,
    WX10841,WX10840,WX10843,WX10842,WX10845,WX10844,WX10847,WX10846,WX10849,
    WX10848,WX10851,WX10850,WX10853,WX10852,WX10855,WX10854,WX10857,WX10856,
    WX10859,WX10858,WX10861,WX10860,WX10863,WX10862,WX10865,WX10864,WX10867,
    WX10866,WX10869,WX10868,WX10871,WX10870,WX10873,WX10872,WX10875,WX10874,
    WX10877,WX10876,WX10879,WX10878,WX10881,WX10880,WX10883,WX10882,WX10885,
    WX10884,WX10887,WX10886,WX10889,WX10888,WX10891,WX10890,WX10989,WX10988,
    WX10991,WX10990,WX10993,WX10992,WX10995,WX10994,WX10997,WX10996,WX10999,
    WX10998,WX11001,WX11000,WX11003,WX11002,WX11005,WX11004,WX11007,WX11006,
    WX11009,WX11008,WX11011,WX11010,WX11013,WX11012,WX11015,WX11014,WX11017,
    WX11016,WX11019,WX11018,WX11021,WX11020,WX11023,WX11022,WX11025,WX11024,
    WX11027,WX11026,WX11029,WX11028,WX11031,WX11030,WX11033,WX11032,WX11035,
    WX11034,WX11037,WX11036,WX11039,WX11038,WX11041,WX11040,WX11043,WX11042,
    WX11045,WX11044,WX11047,WX11046,WX11049,WX11048,WX11051,WX11050,WX11053,
    WX11052,WX11055,WX11054,WX11057,WX11056,WX11059,WX11058,WX11061,WX11060,
    WX11063,WX11062,WX11065,WX11064,WX11067,WX11066,WX11069,WX11068,WX11071,
    WX11070,WX11073,WX11072,WX11075,WX11074,WX11077,WX11076,WX11079,WX11078,
    WX11081,WX11080,WX11083,WX11082,WX11085,WX11084,WX11087,WX11086,WX11089,
    WX11088,WX11091,WX11090,WX11093,WX11092,WX11095,WX11094,WX11097,WX11096,
    WX11099,WX11098,WX11101,WX11100,WX11103,WX11102,WX11105,WX11104,WX11107,
    WX11106,WX11109,WX11108,WX11111,WX11110,WX11113,WX11112,WX11115,WX11114,
    WX11117,WX11116,WX11119,WX11118,WX11121,WX11120,WX11123,WX11122,WX11125,
    WX11124,WX11127,WX11126,WX11129,WX11128,WX11131,WX11130,WX11133,WX11132,
    WX11135,WX11134,WX11137,WX11136,WX11139,WX11138,WX11141,WX11140,WX11143,
    WX11142,WX11145,WX11144,WX11147,WX11146,WX11149,WX11148,WX11151,WX11150,
    WX11153,WX11152,WX11155,WX11154,WX11157,WX11156,WX11159,WX11158,WX11161,
    WX11160,WX11163,WX11162,WX11165,WX11164,WX11167,WX11166,WX11169,WX11168,
    WX11171,WX11170,WX11173,WX11172,WX11175,WX11174,WX11177,WX11176,WX11179,
    WX11178,WX11181,WX11180,WX11183,WX11182,WX11185,WX11184,WX11187,WX11186,
    WX11189,WX11188,WX11191,WX11190,WX11193,WX11192,WX11195,WX11194,WX11197,
    WX11196,WX11199,WX11198,WX11201,WX11200,WX11203,WX11202,WX11205,WX11204,
    WX11207,WX11206,WX11209,WX11208,WX11211,WX11210,WX11213,WX11212,WX11215,
    WX11214,WX11217,WX11216,WX11219,WX11218,WX11221,WX11220,WX11223,WX11222,
    WX11225,WX11224,WX11227,WX11226,WX11229,WX11228,WX11231,WX11230,WX11233,
    WX11232,WX11235,WX11234,WX11237,WX11236,WX11239,WX11238,WX11241,WX11240,
    WX11243,WX11242,WX11608,WX11610,WX11612,WX11614,WX11616,WX11618,WX11620,
    WX11622,WX11624,WX11626,WX11628,WX11630,WX11632,WX11634,WX11636,WX11638,
    WX11640,WX11642,WX11644,WX11646,WX11648,WX11650,WX11652,WX11654,WX11656,
    WX11658,WX11660,WX11662,WX11664,WX11666,WX11668,WX11670,WX37,WX1003,WX41,
    WX1004,WX45,WX47,WX38,WX48,WX51,WX55,WX59,WX61,WX52,WX62,WX65,WX69,WX73,
    WX75,WX66,WX76,WX79,WX83,WX87,WX89,WX80,WX90,WX93,WX97,WX101,WX103,WX94,
    WX104,WX107,WX111,WX115,WX117,WX108,WX118,WX121,WX125,WX129,WX131,WX122,
    WX132,WX135,WX139,WX143,WX145,WX136,WX146,WX149,WX153,WX157,WX159,WX150,
    WX160,WX163,WX167,WX171,WX173,WX164,WX174,WX177,WX181,WX185,WX187,WX178,
    WX188,WX191,WX195,WX199,WX201,WX192,WX202,WX205,WX209,WX213,WX215,WX206,
    WX216,WX219,WX223,WX227,WX229,WX220,WX230,WX233,WX237,WX241,WX243,WX234,
    WX244,WX247,WX251,WX255,WX257,WX248,WX258,WX261,WX265,WX269,WX271,WX262,
    WX272,WX275,WX279,WX283,WX285,WX276,WX286,WX289,WX293,WX297,WX299,WX290,
    WX300,WX303,WX307,WX311,WX313,WX304,WX314,WX317,WX321,WX325,WX327,WX318,
    WX328,WX331,WX335,WX339,WX341,WX332,WX342,WX345,WX349,WX353,WX355,WX346,
    WX356,WX359,WX363,WX367,WX369,WX360,WX370,WX373,WX377,WX381,WX383,WX374,
    WX384,WX387,WX391,WX395,WX397,WX388,WX398,WX401,WX405,WX409,WX411,WX402,
    WX412,WX415,WX419,WX423,WX425,WX416,WX426,WX429,WX433,WX437,WX439,WX430,
    WX440,WX443,WX447,WX451,WX453,WX444,WX454,WX457,WX461,WX465,WX467,WX458,
    WX468,WX471,WX475,WX479,WX481,WX472,WX482,WX483,WX548,WX965,WX549,WX967,
    WX550,WX969,WX551,WX971,WX552,WX973,WX553,WX975,WX554,WX977,WX555,WX979,
    WX556,WX981,WX557,WX983,WX558,WX985,WX559,WX987,WX560,WX989,WX561,WX991,
    WX562,WX993,WX563,WX995,WX564,WX933,WX565,WX935,WX566,WX937,WX567,WX939,
    WX568,WX941,WX569,WX943,WX570,WX945,WX571,WX947,WX572,WX949,WX573,WX951,
    WX574,WX953,WX575,WX955,WX576,WX957,WX577,WX959,WX578,WX961,WX579,WX963,
    WX580,WX581,WX582,WX583,WX584,WX585,WX586,WX587,WX588,WX589,WX590,WX591,
    WX592,WX593,WX594,WX595,WX596,WX597,WX598,WX599,WX600,WX601,WX602,WX603,
    WX604,WX605,WX606,WX607,WX608,WX609,WX610,WX611,WX612,WX613,WX614,WX615,
    WX616,WX617,WX618,WX619,WX620,WX621,WX622,WX623,WX624,WX625,WX626,WX627,
    WX628,WX629,WX630,WX631,WX632,WX633,WX634,WX635,WX636,WX637,WX638,WX639,
    WX640,WX641,WX642,WX643,WX932,WX916,WX934,WX917,WX936,WX918,WX938,WX919,
    WX940,WX920,WX942,WX921,WX944,WX922,WX946,WX923,WX948,WX924,WX950,WX925,
    WX952,WX926,WX954,WX927,WX956,WX928,WX958,WX929,WX960,WX930,WX962,WX931,
    WX964,WX900,WX966,WX901,WX968,WX902,WX970,WX903,WX972,WX904,WX974,WX905,
    WX976,WX906,WX978,WX907,WX980,WX908,WX982,WX909,WX984,WX910,WX986,WX911,
    WX988,WX912,WX990,WX913,WX992,WX914,WX994,WX915,WX996,WX997,WX998,WX999,
    WX1000,WX1001,WX1002,WX1005,WX1009,WX1011,WX1010,WX1016,WX1018,WX1017,
    WX1023,WX1025,WX1024,WX1030,WX1032,WX1031,WX1037,WX1039,WX1038,WX1044,
    WX1046,WX1045,WX1051,WX1053,WX1052,WX1058,WX1060,WX1059,WX1065,WX1067,
    WX1066,WX1072,WX1074,WX1073,WX1079,WX1081,WX1080,WX1086,WX1088,WX1087,
    WX1093,WX1095,WX1094,WX1100,WX1102,WX1101,WX1107,WX1109,WX1108,WX1114,
    WX1116,WX1115,WX1121,WX1123,WX1122,WX1128,WX1130,WX1129,WX1135,WX1137,
    WX1136,WX1142,WX1144,WX1143,WX1149,WX1151,WX1150,WX1156,WX1158,WX1157,
    WX1163,WX1165,WX1164,WX1170,WX1172,WX1171,WX1177,WX1179,WX1178,WX1184,
    WX1186,WX1185,WX1191,WX1193,WX1192,WX1198,WX1200,WX1199,WX1205,WX1207,
    WX1206,WX1212,WX1214,WX1213,WX1219,WX1221,WX1220,WX1226,WX1228,WX1227,
    WX1230,WX1263,WX1330,WX2296,WX1334,WX2297,WX1338,WX1340,WX1331,WX1341,
    WX1344,WX1348,WX1352,WX1354,WX1345,WX1355,WX1358,WX1362,WX1366,WX1368,
    WX1359,WX1369,WX1372,WX1376,WX1380,WX1382,WX1373,WX1383,WX1386,WX1390,
    WX1394,WX1396,WX1387,WX1397,WX1400,WX1404,WX1408,WX1410,WX1401,WX1411,
    WX1414,WX1418,WX1422,WX1424,WX1415,WX1425,WX1428,WX1432,WX1436,WX1438,
    WX1429,WX1439,WX1442,WX1446,WX1450,WX1452,WX1443,WX1453,WX1456,WX1460,
    WX1464,WX1466,WX1457,WX1467,WX1470,WX1474,WX1478,WX1480,WX1471,WX1481,
    WX1484,WX1488,WX1492,WX1494,WX1485,WX1495,WX1498,WX1502,WX1506,WX1508,
    WX1499,WX1509,WX1512,WX1516,WX1520,WX1522,WX1513,WX1523,WX1526,WX1530,
    WX1534,WX1536,WX1527,WX1537,WX1540,WX1544,WX1548,WX1550,WX1541,WX1551,
    WX1554,WX1558,WX1562,WX1564,WX1555,WX1565,WX1568,WX1572,WX1576,WX1578,
    WX1569,WX1579,WX1582,WX1586,WX1590,WX1592,WX1583,WX1593,WX1596,WX1600,
    WX1604,WX1606,WX1597,WX1607,WX1610,WX1614,WX1618,WX1620,WX1611,WX1621,
    WX1624,WX1628,WX1632,WX1634,WX1625,WX1635,WX1638,WX1642,WX1646,WX1648,
    WX1639,WX1649,WX1652,WX1656,WX1660,WX1662,WX1653,WX1663,WX1666,WX1670,
    WX1674,WX1676,WX1667,WX1677,WX1680,WX1684,WX1688,WX1690,WX1681,WX1691,
    WX1694,WX1698,WX1702,WX1704,WX1695,WX1705,WX1708,WX1712,WX1716,WX1718,
    WX1709,WX1719,WX1722,WX1726,WX1730,WX1732,WX1723,WX1733,WX1736,WX1740,
    WX1744,WX1746,WX1737,WX1747,WX1750,WX1754,WX1758,WX1760,WX1751,WX1761,
    WX1764,WX1768,WX1772,WX1774,WX1765,WX1775,WX1776,WX1841,WX2258,WX1842,
    WX2260,WX1843,WX2262,WX1844,WX2264,WX1845,WX2266,WX1846,WX2268,WX1847,
    WX2270,WX1848,WX2272,WX1849,WX2274,WX1850,WX2276,WX1851,WX2278,WX1852,
    WX2280,WX1853,WX2282,WX1854,WX2284,WX1855,WX2286,WX1856,WX2288,WX1857,
    WX2226,WX1858,WX2228,WX1859,WX2230,WX1860,WX2232,WX1861,WX2234,WX1862,
    WX2236,WX1863,WX2238,WX1864,WX2240,WX1865,WX2242,WX1866,WX2244,WX1867,
    WX2246,WX1868,WX2248,WX1869,WX2250,WX1870,WX2252,WX1871,WX2254,WX1872,
    WX2256,WX1873,WX1874,WX1875,WX1876,WX1877,WX1878,WX1879,WX1880,WX1881,
    WX1882,WX1883,WX1884,WX1885,WX1886,WX1887,WX1888,WX1889,WX1890,WX1891,
    WX1892,WX1893,WX1894,WX1895,WX1896,WX1897,WX1898,WX1899,WX1900,WX1901,
    WX1902,WX1903,WX1904,WX1905,WX1906,WX1907,WX1908,WX1909,WX1910,WX1911,
    WX1912,WX1913,WX1914,WX1915,WX1916,WX1917,WX1918,WX1919,WX1920,WX1921,
    WX1922,WX1923,WX1924,WX1925,WX1926,WX1927,WX1928,WX1929,WX1930,WX1931,
    WX1932,WX1933,WX1934,WX1935,WX1936,WX2225,WX2209,WX2227,WX2210,WX2229,
    WX2211,WX2231,WX2212,WX2233,WX2213,WX2235,WX2214,WX2237,WX2215,WX2239,
    WX2216,WX2241,WX2217,WX2243,WX2218,WX2245,WX2219,WX2247,WX2220,WX2249,
    WX2221,WX2251,WX2222,WX2253,WX2223,WX2255,WX2224,WX2257,WX2193,WX2259,
    WX2194,WX2261,WX2195,WX2263,WX2196,WX2265,WX2197,WX2267,WX2198,WX2269,
    WX2199,WX2271,WX2200,WX2273,WX2201,WX2275,WX2202,WX2277,WX2203,WX2279,
    WX2204,WX2281,WX2205,WX2283,WX2206,WX2285,WX2207,WX2287,WX2208,WX2289,
    WX2290,WX2291,WX2292,WX2293,WX2294,WX2295,WX2298,WX2302,WX2304,WX2303,
    WX2305,WX2309,WX2311,WX2310,WX2312,WX2316,WX2318,WX2317,WX2319,WX2323,
    WX2325,WX2324,WX2326,WX2330,WX2332,WX2331,WX2333,WX2337,WX2339,WX2338,
    WX2340,WX2344,WX2346,WX2345,WX2347,WX2351,WX2353,WX2352,WX2354,WX2358,
    WX2360,WX2359,WX2361,WX2365,WX2367,WX2366,WX2368,WX2372,WX2374,WX2373,
    WX2375,WX2379,WX2381,WX2380,WX2382,WX2386,WX2388,WX2387,WX2389,WX2393,
    WX2395,WX2394,WX2396,WX2400,WX2402,WX2401,WX2403,WX2407,WX2409,WX2408,
    WX2410,WX2414,WX2416,WX2415,WX2417,WX2421,WX2423,WX2422,WX2424,WX2428,
    WX2430,WX2429,WX2431,WX2435,WX2437,WX2436,WX2438,WX2442,WX2444,WX2443,
    WX2445,WX2449,WX2451,WX2450,WX2452,WX2456,WX2458,WX2457,WX2459,WX2463,
    WX2465,WX2464,WX2466,WX2470,WX2472,WX2471,WX2473,WX2477,WX2479,WX2478,
    WX2480,WX2484,WX2486,WX2485,WX2487,WX2491,WX2493,WX2492,WX2494,WX2498,
    WX2500,WX2499,WX2501,WX2505,WX2507,WX2506,WX2508,WX2512,WX2514,WX2513,
    WX2515,WX2519,WX2521,WX2520,WX2522,WX2523,WX2556,WX2623,WX3589,WX2627,
    WX3590,WX2631,WX2633,WX2624,WX2634,WX2637,WX2641,WX2645,WX2647,WX2638,
    WX2648,WX2651,WX2655,WX2659,WX2661,WX2652,WX2662,WX2665,WX2669,WX2673,
    WX2675,WX2666,WX2676,WX2679,WX2683,WX2687,WX2689,WX2680,WX2690,WX2693,
    WX2697,WX2701,WX2703,WX2694,WX2704,WX2707,WX2711,WX2715,WX2717,WX2708,
    WX2718,WX2721,WX2725,WX2729,WX2731,WX2722,WX2732,WX2735,WX2739,WX2743,
    WX2745,WX2736,WX2746,WX2749,WX2753,WX2757,WX2759,WX2750,WX2760,WX2763,
    WX2767,WX2771,WX2773,WX2764,WX2774,WX2777,WX2781,WX2785,WX2787,WX2778,
    WX2788,WX2791,WX2795,WX2799,WX2801,WX2792,WX2802,WX2805,WX2809,WX2813,
    WX2815,WX2806,WX2816,WX2819,WX2823,WX2827,WX2829,WX2820,WX2830,WX2833,
    WX2837,WX2841,WX2843,WX2834,WX2844,WX2847,WX2851,WX2855,WX2857,WX2848,
    WX2858,WX2861,WX2865,WX2869,WX2871,WX2862,WX2872,WX2875,WX2879,WX2883,
    WX2885,WX2876,WX2886,WX2889,WX2893,WX2897,WX2899,WX2890,WX2900,WX2903,
    WX2907,WX2911,WX2913,WX2904,WX2914,WX2917,WX2921,WX2925,WX2927,WX2918,
    WX2928,WX2931,WX2935,WX2939,WX2941,WX2932,WX2942,WX2945,WX2949,WX2953,
    WX2955,WX2946,WX2956,WX2959,WX2963,WX2967,WX2969,WX2960,WX2970,WX2973,
    WX2977,WX2981,WX2983,WX2974,WX2984,WX2987,WX2991,WX2995,WX2997,WX2988,
    WX2998,WX3001,WX3005,WX3009,WX3011,WX3002,WX3012,WX3015,WX3019,WX3023,
    WX3025,WX3016,WX3026,WX3029,WX3033,WX3037,WX3039,WX3030,WX3040,WX3043,
    WX3047,WX3051,WX3053,WX3044,WX3054,WX3057,WX3061,WX3065,WX3067,WX3058,
    WX3068,WX3069,WX3134,WX3551,WX3135,WX3553,WX3136,WX3555,WX3137,WX3557,
    WX3138,WX3559,WX3139,WX3561,WX3140,WX3563,WX3141,WX3565,WX3142,WX3567,
    WX3143,WX3569,WX3144,WX3571,WX3145,WX3573,WX3146,WX3575,WX3147,WX3577,
    WX3148,WX3579,WX3149,WX3581,WX3150,WX3519,WX3151,WX3521,WX3152,WX3523,
    WX3153,WX3525,WX3154,WX3527,WX3155,WX3529,WX3156,WX3531,WX3157,WX3533,
    WX3158,WX3535,WX3159,WX3537,WX3160,WX3539,WX3161,WX3541,WX3162,WX3543,
    WX3163,WX3545,WX3164,WX3547,WX3165,WX3549,WX3166,WX3167,WX3168,WX3169,
    WX3170,WX3171,WX3172,WX3173,WX3174,WX3175,WX3176,WX3177,WX3178,WX3179,
    WX3180,WX3181,WX3182,WX3183,WX3184,WX3185,WX3186,WX3187,WX3188,WX3189,
    WX3190,WX3191,WX3192,WX3193,WX3194,WX3195,WX3196,WX3197,WX3198,WX3199,
    WX3200,WX3201,WX3202,WX3203,WX3204,WX3205,WX3206,WX3207,WX3208,WX3209,
    WX3210,WX3211,WX3212,WX3213,WX3214,WX3215,WX3216,WX3217,WX3218,WX3219,
    WX3220,WX3221,WX3222,WX3223,WX3224,WX3225,WX3226,WX3227,WX3228,WX3229,
    WX3518,WX3502,WX3520,WX3503,WX3522,WX3504,WX3524,WX3505,WX3526,WX3506,
    WX3528,WX3507,WX3530,WX3508,WX3532,WX3509,WX3534,WX3510,WX3536,WX3511,
    WX3538,WX3512,WX3540,WX3513,WX3542,WX3514,WX3544,WX3515,WX3546,WX3516,
    WX3548,WX3517,WX3550,WX3486,WX3552,WX3487,WX3554,WX3488,WX3556,WX3489,
    WX3558,WX3490,WX3560,WX3491,WX3562,WX3492,WX3564,WX3493,WX3566,WX3494,
    WX3568,WX3495,WX3570,WX3496,WX3572,WX3497,WX3574,WX3498,WX3576,WX3499,
    WX3578,WX3500,WX3580,WX3501,WX3582,WX3583,WX3584,WX3585,WX3586,WX3587,
    WX3588,WX3591,WX3595,WX3597,WX3596,WX3598,WX3602,WX3604,WX3603,WX3605,
    WX3609,WX3611,WX3610,WX3612,WX3616,WX3618,WX3617,WX3619,WX3623,WX3625,
    WX3624,WX3626,WX3630,WX3632,WX3631,WX3633,WX3637,WX3639,WX3638,WX3640,
    WX3644,WX3646,WX3645,WX3647,WX3651,WX3653,WX3652,WX3654,WX3658,WX3660,
    WX3659,WX3661,WX3665,WX3667,WX3666,WX3668,WX3672,WX3674,WX3673,WX3675,
    WX3679,WX3681,WX3680,WX3682,WX3686,WX3688,WX3687,WX3689,WX3693,WX3695,
    WX3694,WX3696,WX3700,WX3702,WX3701,WX3703,WX3707,WX3709,WX3708,WX3710,
    WX3714,WX3716,WX3715,WX3717,WX3721,WX3723,WX3722,WX3724,WX3728,WX3730,
    WX3729,WX3731,WX3735,WX3737,WX3736,WX3738,WX3742,WX3744,WX3743,WX3745,
    WX3749,WX3751,WX3750,WX3752,WX3756,WX3758,WX3757,WX3759,WX3763,WX3765,
    WX3764,WX3766,WX3770,WX3772,WX3771,WX3773,WX3777,WX3779,WX3778,WX3780,
    WX3784,WX3786,WX3785,WX3787,WX3791,WX3793,WX3792,WX3794,WX3798,WX3800,
    WX3799,WX3801,WX3805,WX3807,WX3806,WX3808,WX3812,WX3814,WX3813,WX3815,
    WX3816,WX3849,WX3916,WX4882,WX3920,WX4883,WX3924,WX3926,WX3917,WX3927,
    WX3930,WX3934,WX3938,WX3940,WX3931,WX3941,WX3944,WX3948,WX3952,WX3954,
    WX3945,WX3955,WX3958,WX3962,WX3966,WX3968,WX3959,WX3969,WX3972,WX3976,
    WX3980,WX3982,WX3973,WX3983,WX3986,WX3990,WX3994,WX3996,WX3987,WX3997,
    WX4000,WX4004,WX4008,WX4010,WX4001,WX4011,WX4014,WX4018,WX4022,WX4024,
    WX4015,WX4025,WX4028,WX4032,WX4036,WX4038,WX4029,WX4039,WX4042,WX4046,
    WX4050,WX4052,WX4043,WX4053,WX4056,WX4060,WX4064,WX4066,WX4057,WX4067,
    WX4070,WX4074,WX4078,WX4080,WX4071,WX4081,WX4084,WX4088,WX4092,WX4094,
    WX4085,WX4095,WX4098,WX4102,WX4106,WX4108,WX4099,WX4109,WX4112,WX4116,
    WX4120,WX4122,WX4113,WX4123,WX4126,WX4130,WX4134,WX4136,WX4127,WX4137,
    WX4140,WX4144,WX4148,WX4150,WX4141,WX4151,WX4154,WX4158,WX4162,WX4164,
    WX4155,WX4165,WX4168,WX4172,WX4176,WX4178,WX4169,WX4179,WX4182,WX4186,
    WX4190,WX4192,WX4183,WX4193,WX4196,WX4200,WX4204,WX4206,WX4197,WX4207,
    WX4210,WX4214,WX4218,WX4220,WX4211,WX4221,WX4224,WX4228,WX4232,WX4234,
    WX4225,WX4235,WX4238,WX4242,WX4246,WX4248,WX4239,WX4249,WX4252,WX4256,
    WX4260,WX4262,WX4253,WX4263,WX4266,WX4270,WX4274,WX4276,WX4267,WX4277,
    WX4280,WX4284,WX4288,WX4290,WX4281,WX4291,WX4294,WX4298,WX4302,WX4304,
    WX4295,WX4305,WX4308,WX4312,WX4316,WX4318,WX4309,WX4319,WX4322,WX4326,
    WX4330,WX4332,WX4323,WX4333,WX4336,WX4340,WX4344,WX4346,WX4337,WX4347,
    WX4350,WX4354,WX4358,WX4360,WX4351,WX4361,WX4362,WX4427,WX4844,WX4428,
    WX4846,WX4429,WX4848,WX4430,WX4850,WX4431,WX4852,WX4432,WX4854,WX4433,
    WX4856,WX4434,WX4858,WX4435,WX4860,WX4436,WX4862,WX4437,WX4864,WX4438,
    WX4866,WX4439,WX4868,WX4440,WX4870,WX4441,WX4872,WX4442,WX4874,WX4443,
    WX4812,WX4444,WX4814,WX4445,WX4816,WX4446,WX4818,WX4447,WX4820,WX4448,
    WX4822,WX4449,WX4824,WX4450,WX4826,WX4451,WX4828,WX4452,WX4830,WX4453,
    WX4832,WX4454,WX4834,WX4455,WX4836,WX4456,WX4838,WX4457,WX4840,WX4458,
    WX4842,WX4459,WX4460,WX4461,WX4462,WX4463,WX4464,WX4465,WX4466,WX4467,
    WX4468,WX4469,WX4470,WX4471,WX4472,WX4473,WX4474,WX4475,WX4476,WX4477,
    WX4478,WX4479,WX4480,WX4481,WX4482,WX4483,WX4484,WX4485,WX4486,WX4487,
    WX4488,WX4489,WX4490,WX4491,WX4492,WX4493,WX4494,WX4495,WX4496,WX4497,
    WX4498,WX4499,WX4500,WX4501,WX4502,WX4503,WX4504,WX4505,WX4506,WX4507,
    WX4508,WX4509,WX4510,WX4511,WX4512,WX4513,WX4514,WX4515,WX4516,WX4517,
    WX4518,WX4519,WX4520,WX4521,WX4522,WX4811,WX4795,WX4813,WX4796,WX4815,
    WX4797,WX4817,WX4798,WX4819,WX4799,WX4821,WX4800,WX4823,WX4801,WX4825,
    WX4802,WX4827,WX4803,WX4829,WX4804,WX4831,WX4805,WX4833,WX4806,WX4835,
    WX4807,WX4837,WX4808,WX4839,WX4809,WX4841,WX4810,WX4843,WX4779,WX4845,
    WX4780,WX4847,WX4781,WX4849,WX4782,WX4851,WX4783,WX4853,WX4784,WX4855,
    WX4785,WX4857,WX4786,WX4859,WX4787,WX4861,WX4788,WX4863,WX4789,WX4865,
    WX4790,WX4867,WX4791,WX4869,WX4792,WX4871,WX4793,WX4873,WX4794,WX4875,
    WX4876,WX4877,WX4878,WX4879,WX4880,WX4881,WX4884,WX4888,WX4890,WX4889,
    WX4891,WX4895,WX4897,WX4896,WX4898,WX4902,WX4904,WX4903,WX4905,WX4909,
    WX4911,WX4910,WX4912,WX4916,WX4918,WX4917,WX4919,WX4923,WX4925,WX4924,
    WX4926,WX4930,WX4932,WX4931,WX4933,WX4937,WX4939,WX4938,WX4940,WX4944,
    WX4946,WX4945,WX4947,WX4951,WX4953,WX4952,WX4954,WX4958,WX4960,WX4959,
    WX4961,WX4965,WX4967,WX4966,WX4968,WX4972,WX4974,WX4973,WX4975,WX4979,
    WX4981,WX4980,WX4982,WX4986,WX4988,WX4987,WX4989,WX4993,WX4995,WX4994,
    WX4996,WX5000,WX5002,WX5001,WX5003,WX5007,WX5009,WX5008,WX5010,WX5014,
    WX5016,WX5015,WX5017,WX5021,WX5023,WX5022,WX5024,WX5028,WX5030,WX5029,
    WX5031,WX5035,WX5037,WX5036,WX5038,WX5042,WX5044,WX5043,WX5045,WX5049,
    WX5051,WX5050,WX5052,WX5056,WX5058,WX5057,WX5059,WX5063,WX5065,WX5064,
    WX5066,WX5070,WX5072,WX5071,WX5073,WX5077,WX5079,WX5078,WX5080,WX5084,
    WX5086,WX5085,WX5087,WX5091,WX5093,WX5092,WX5094,WX5098,WX5100,WX5099,
    WX5101,WX5105,WX5107,WX5106,WX5108,WX5109,WX5142,WX5209,WX6175,WX5213,
    WX6176,WX5217,WX5219,WX5210,WX5220,WX5223,WX5227,WX5231,WX5233,WX5224,
    WX5234,WX5237,WX5241,WX5245,WX5247,WX5238,WX5248,WX5251,WX5255,WX5259,
    WX5261,WX5252,WX5262,WX5265,WX5269,WX5273,WX5275,WX5266,WX5276,WX5279,
    WX5283,WX5287,WX5289,WX5280,WX5290,WX5293,WX5297,WX5301,WX5303,WX5294,
    WX5304,WX5307,WX5311,WX5315,WX5317,WX5308,WX5318,WX5321,WX5325,WX5329,
    WX5331,WX5322,WX5332,WX5335,WX5339,WX5343,WX5345,WX5336,WX5346,WX5349,
    WX5353,WX5357,WX5359,WX5350,WX5360,WX5363,WX5367,WX5371,WX5373,WX5364,
    WX5374,WX5377,WX5381,WX5385,WX5387,WX5378,WX5388,WX5391,WX5395,WX5399,
    WX5401,WX5392,WX5402,WX5405,WX5409,WX5413,WX5415,WX5406,WX5416,WX5419,
    WX5423,WX5427,WX5429,WX5420,WX5430,WX5433,WX5437,WX5441,WX5443,WX5434,
    WX5444,WX5447,WX5451,WX5455,WX5457,WX5448,WX5458,WX5461,WX5465,WX5469,
    WX5471,WX5462,WX5472,WX5475,WX5479,WX5483,WX5485,WX5476,WX5486,WX5489,
    WX5493,WX5497,WX5499,WX5490,WX5500,WX5503,WX5507,WX5511,WX5513,WX5504,
    WX5514,WX5517,WX5521,WX5525,WX5527,WX5518,WX5528,WX5531,WX5535,WX5539,
    WX5541,WX5532,WX5542,WX5545,WX5549,WX5553,WX5555,WX5546,WX5556,WX5559,
    WX5563,WX5567,WX5569,WX5560,WX5570,WX5573,WX5577,WX5581,WX5583,WX5574,
    WX5584,WX5587,WX5591,WX5595,WX5597,WX5588,WX5598,WX5601,WX5605,WX5609,
    WX5611,WX5602,WX5612,WX5615,WX5619,WX5623,WX5625,WX5616,WX5626,WX5629,
    WX5633,WX5637,WX5639,WX5630,WX5640,WX5643,WX5647,WX5651,WX5653,WX5644,
    WX5654,WX5655,WX5720,WX6137,WX5721,WX6139,WX5722,WX6141,WX5723,WX6143,
    WX5724,WX6145,WX5725,WX6147,WX5726,WX6149,WX5727,WX6151,WX5728,WX6153,
    WX5729,WX6155,WX5730,WX6157,WX5731,WX6159,WX5732,WX6161,WX5733,WX6163,
    WX5734,WX6165,WX5735,WX6167,WX5736,WX6105,WX5737,WX6107,WX5738,WX6109,
    WX5739,WX6111,WX5740,WX6113,WX5741,WX6115,WX5742,WX6117,WX5743,WX6119,
    WX5744,WX6121,WX5745,WX6123,WX5746,WX6125,WX5747,WX6127,WX5748,WX6129,
    WX5749,WX6131,WX5750,WX6133,WX5751,WX6135,WX5752,WX5753,WX5754,WX5755,
    WX5756,WX5757,WX5758,WX5759,WX5760,WX5761,WX5762,WX5763,WX5764,WX5765,
    WX5766,WX5767,WX5768,WX5769,WX5770,WX5771,WX5772,WX5773,WX5774,WX5775,
    WX5776,WX5777,WX5778,WX5779,WX5780,WX5781,WX5782,WX5783,WX5784,WX5785,
    WX5786,WX5787,WX5788,WX5789,WX5790,WX5791,WX5792,WX5793,WX5794,WX5795,
    WX5796,WX5797,WX5798,WX5799,WX5800,WX5801,WX5802,WX5803,WX5804,WX5805,
    WX5806,WX5807,WX5808,WX5809,WX5810,WX5811,WX5812,WX5813,WX5814,WX5815,
    WX6104,WX6088,WX6106,WX6089,WX6108,WX6090,WX6110,WX6091,WX6112,WX6092,
    WX6114,WX6093,WX6116,WX6094,WX6118,WX6095,WX6120,WX6096,WX6122,WX6097,
    WX6124,WX6098,WX6126,WX6099,WX6128,WX6100,WX6130,WX6101,WX6132,WX6102,
    WX6134,WX6103,WX6136,WX6072,WX6138,WX6073,WX6140,WX6074,WX6142,WX6075,
    WX6144,WX6076,WX6146,WX6077,WX6148,WX6078,WX6150,WX6079,WX6152,WX6080,
    WX6154,WX6081,WX6156,WX6082,WX6158,WX6083,WX6160,WX6084,WX6162,WX6085,
    WX6164,WX6086,WX6166,WX6087,WX6168,WX6169,WX6170,WX6171,WX6172,WX6173,
    WX6174,WX6177,WX6181,WX6183,WX6182,WX6184,WX6188,WX6190,WX6189,WX6191,
    WX6195,WX6197,WX6196,WX6198,WX6202,WX6204,WX6203,WX6205,WX6209,WX6211,
    WX6210,WX6212,WX6216,WX6218,WX6217,WX6219,WX6223,WX6225,WX6224,WX6226,
    WX6230,WX6232,WX6231,WX6233,WX6237,WX6239,WX6238,WX6240,WX6244,WX6246,
    WX6245,WX6247,WX6251,WX6253,WX6252,WX6254,WX6258,WX6260,WX6259,WX6261,
    WX6265,WX6267,WX6266,WX6268,WX6272,WX6274,WX6273,WX6275,WX6279,WX6281,
    WX6280,WX6282,WX6286,WX6288,WX6287,WX6289,WX6293,WX6295,WX6294,WX6296,
    WX6300,WX6302,WX6301,WX6303,WX6307,WX6309,WX6308,WX6310,WX6314,WX6316,
    WX6315,WX6317,WX6321,WX6323,WX6322,WX6324,WX6328,WX6330,WX6329,WX6331,
    WX6335,WX6337,WX6336,WX6338,WX6342,WX6344,WX6343,WX6345,WX6349,WX6351,
    WX6350,WX6352,WX6356,WX6358,WX6357,WX6359,WX6363,WX6365,WX6364,WX6366,
    WX6370,WX6372,WX6371,WX6373,WX6377,WX6379,WX6378,WX6380,WX6384,WX6386,
    WX6385,WX6387,WX6391,WX6393,WX6392,WX6394,WX6398,WX6400,WX6399,WX6401,
    WX6402,WX6435,WX6502,WX7468,WX6506,WX7469,WX6510,WX6512,WX6503,WX6513,
    WX6516,WX6520,WX6524,WX6526,WX6517,WX6527,WX6530,WX6534,WX6538,WX6540,
    WX6531,WX6541,WX6544,WX6548,WX6552,WX6554,WX6545,WX6555,WX6558,WX6562,
    WX6566,WX6568,WX6559,WX6569,WX6572,WX6576,WX6580,WX6582,WX6573,WX6583,
    WX6586,WX6590,WX6594,WX6596,WX6587,WX6597,WX6600,WX6604,WX6608,WX6610,
    WX6601,WX6611,WX6614,WX6618,WX6622,WX6624,WX6615,WX6625,WX6628,WX6632,
    WX6636,WX6638,WX6629,WX6639,WX6642,WX6646,WX6650,WX6652,WX6643,WX6653,
    WX6656,WX6660,WX6664,WX6666,WX6657,WX6667,WX6670,WX6674,WX6678,WX6680,
    WX6671,WX6681,WX6684,WX6688,WX6692,WX6694,WX6685,WX6695,WX6698,WX6702,
    WX6706,WX6708,WX6699,WX6709,WX6712,WX6716,WX6720,WX6722,WX6713,WX6723,
    WX6726,WX6730,WX6734,WX6736,WX6727,WX6737,WX6740,WX6744,WX6748,WX6750,
    WX6741,WX6751,WX6754,WX6758,WX6762,WX6764,WX6755,WX6765,WX6768,WX6772,
    WX6776,WX6778,WX6769,WX6779,WX6782,WX6786,WX6790,WX6792,WX6783,WX6793,
    WX6796,WX6800,WX6804,WX6806,WX6797,WX6807,WX6810,WX6814,WX6818,WX6820,
    WX6811,WX6821,WX6824,WX6828,WX6832,WX6834,WX6825,WX6835,WX6838,WX6842,
    WX6846,WX6848,WX6839,WX6849,WX6852,WX6856,WX6860,WX6862,WX6853,WX6863,
    WX6866,WX6870,WX6874,WX6876,WX6867,WX6877,WX6880,WX6884,WX6888,WX6890,
    WX6881,WX6891,WX6894,WX6898,WX6902,WX6904,WX6895,WX6905,WX6908,WX6912,
    WX6916,WX6918,WX6909,WX6919,WX6922,WX6926,WX6930,WX6932,WX6923,WX6933,
    WX6936,WX6940,WX6944,WX6946,WX6937,WX6947,WX6948,WX7013,WX7430,WX7014,
    WX7432,WX7015,WX7434,WX7016,WX7436,WX7017,WX7438,WX7018,WX7440,WX7019,
    WX7442,WX7020,WX7444,WX7021,WX7446,WX7022,WX7448,WX7023,WX7450,WX7024,
    WX7452,WX7025,WX7454,WX7026,WX7456,WX7027,WX7458,WX7028,WX7460,WX7029,
    WX7398,WX7030,WX7400,WX7031,WX7402,WX7032,WX7404,WX7033,WX7406,WX7034,
    WX7408,WX7035,WX7410,WX7036,WX7412,WX7037,WX7414,WX7038,WX7416,WX7039,
    WX7418,WX7040,WX7420,WX7041,WX7422,WX7042,WX7424,WX7043,WX7426,WX7044,
    WX7428,WX7045,WX7046,WX7047,WX7048,WX7049,WX7050,WX7051,WX7052,WX7053,
    WX7054,WX7055,WX7056,WX7057,WX7058,WX7059,WX7060,WX7061,WX7062,WX7063,
    WX7064,WX7065,WX7066,WX7067,WX7068,WX7069,WX7070,WX7071,WX7072,WX7073,
    WX7074,WX7075,WX7076,WX7077,WX7078,WX7079,WX7080,WX7081,WX7082,WX7083,
    WX7084,WX7085,WX7086,WX7087,WX7088,WX7089,WX7090,WX7091,WX7092,WX7093,
    WX7094,WX7095,WX7096,WX7097,WX7098,WX7099,WX7100,WX7101,WX7102,WX7103,
    WX7104,WX7105,WX7106,WX7107,WX7108,WX7397,WX7381,WX7399,WX7382,WX7401,
    WX7383,WX7403,WX7384,WX7405,WX7385,WX7407,WX7386,WX7409,WX7387,WX7411,
    WX7388,WX7413,WX7389,WX7415,WX7390,WX7417,WX7391,WX7419,WX7392,WX7421,
    WX7393,WX7423,WX7394,WX7425,WX7395,WX7427,WX7396,WX7429,WX7365,WX7431,
    WX7366,WX7433,WX7367,WX7435,WX7368,WX7437,WX7369,WX7439,WX7370,WX7441,
    WX7371,WX7443,WX7372,WX7445,WX7373,WX7447,WX7374,WX7449,WX7375,WX7451,
    WX7376,WX7453,WX7377,WX7455,WX7378,WX7457,WX7379,WX7459,WX7380,WX7461,
    WX7462,WX7463,WX7464,WX7465,WX7466,WX7467,WX7470,WX7474,WX7476,WX7475,
    WX7477,WX7481,WX7483,WX7482,WX7484,WX7488,WX7490,WX7489,WX7491,WX7495,
    WX7497,WX7496,WX7498,WX7502,WX7504,WX7503,WX7505,WX7509,WX7511,WX7510,
    WX7512,WX7516,WX7518,WX7517,WX7519,WX7523,WX7525,WX7524,WX7526,WX7530,
    WX7532,WX7531,WX7533,WX7537,WX7539,WX7538,WX7540,WX7544,WX7546,WX7545,
    WX7547,WX7551,WX7553,WX7552,WX7554,WX7558,WX7560,WX7559,WX7561,WX7565,
    WX7567,WX7566,WX7568,WX7572,WX7574,WX7573,WX7575,WX7579,WX7581,WX7580,
    WX7582,WX7586,WX7588,WX7587,WX7589,WX7593,WX7595,WX7594,WX7596,WX7600,
    WX7602,WX7601,WX7603,WX7607,WX7609,WX7608,WX7610,WX7614,WX7616,WX7615,
    WX7617,WX7621,WX7623,WX7622,WX7624,WX7628,WX7630,WX7629,WX7631,WX7635,
    WX7637,WX7636,WX7638,WX7642,WX7644,WX7643,WX7645,WX7649,WX7651,WX7650,
    WX7652,WX7656,WX7658,WX7657,WX7659,WX7663,WX7665,WX7664,WX7666,WX7670,
    WX7672,WX7671,WX7673,WX7677,WX7679,WX7678,WX7680,WX7684,WX7686,WX7685,
    WX7687,WX7691,WX7693,WX7692,WX7694,WX7695,WX7728,WX7795,WX8761,WX7799,
    WX8762,WX7803,WX7805,WX7796,WX7806,WX7809,WX7813,WX7817,WX7819,WX7810,
    WX7820,WX7823,WX7827,WX7831,WX7833,WX7824,WX7834,WX7837,WX7841,WX7845,
    WX7847,WX7838,WX7848,WX7851,WX7855,WX7859,WX7861,WX7852,WX7862,WX7865,
    WX7869,WX7873,WX7875,WX7866,WX7876,WX7879,WX7883,WX7887,WX7889,WX7880,
    WX7890,WX7893,WX7897,WX7901,WX7903,WX7894,WX7904,WX7907,WX7911,WX7915,
    WX7917,WX7908,WX7918,WX7921,WX7925,WX7929,WX7931,WX7922,WX7932,WX7935,
    WX7939,WX7943,WX7945,WX7936,WX7946,WX7949,WX7953,WX7957,WX7959,WX7950,
    WX7960,WX7963,WX7967,WX7971,WX7973,WX7964,WX7974,WX7977,WX7981,WX7985,
    WX7987,WX7978,WX7988,WX7991,WX7995,WX7999,WX8001,WX7992,WX8002,WX8005,
    WX8009,WX8013,WX8015,WX8006,WX8016,WX8019,WX8023,WX8027,WX8029,WX8020,
    WX8030,WX8033,WX8037,WX8041,WX8043,WX8034,WX8044,WX8047,WX8051,WX8055,
    WX8057,WX8048,WX8058,WX8061,WX8065,WX8069,WX8071,WX8062,WX8072,WX8075,
    WX8079,WX8083,WX8085,WX8076,WX8086,WX8089,WX8093,WX8097,WX8099,WX8090,
    WX8100,WX8103,WX8107,WX8111,WX8113,WX8104,WX8114,WX8117,WX8121,WX8125,
    WX8127,WX8118,WX8128,WX8131,WX8135,WX8139,WX8141,WX8132,WX8142,WX8145,
    WX8149,WX8153,WX8155,WX8146,WX8156,WX8159,WX8163,WX8167,WX8169,WX8160,
    WX8170,WX8173,WX8177,WX8181,WX8183,WX8174,WX8184,WX8187,WX8191,WX8195,
    WX8197,WX8188,WX8198,WX8201,WX8205,WX8209,WX8211,WX8202,WX8212,WX8215,
    WX8219,WX8223,WX8225,WX8216,WX8226,WX8229,WX8233,WX8237,WX8239,WX8230,
    WX8240,WX8241,WX8306,WX8723,WX8307,WX8725,WX8308,WX8727,WX8309,WX8729,
    WX8310,WX8731,WX8311,WX8733,WX8312,WX8735,WX8313,WX8737,WX8314,WX8739,
    WX8315,WX8741,WX8316,WX8743,WX8317,WX8745,WX8318,WX8747,WX8319,WX8749,
    WX8320,WX8751,WX8321,WX8753,WX8322,WX8691,WX8323,WX8693,WX8324,WX8695,
    WX8325,WX8697,WX8326,WX8699,WX8327,WX8701,WX8328,WX8703,WX8329,WX8705,
    WX8330,WX8707,WX8331,WX8709,WX8332,WX8711,WX8333,WX8713,WX8334,WX8715,
    WX8335,WX8717,WX8336,WX8719,WX8337,WX8721,WX8338,WX8339,WX8340,WX8341,
    WX8342,WX8343,WX8344,WX8345,WX8346,WX8347,WX8348,WX8349,WX8350,WX8351,
    WX8352,WX8353,WX8354,WX8355,WX8356,WX8357,WX8358,WX8359,WX8360,WX8361,
    WX8362,WX8363,WX8364,WX8365,WX8366,WX8367,WX8368,WX8369,WX8370,WX8371,
    WX8372,WX8373,WX8374,WX8375,WX8376,WX8377,WX8378,WX8379,WX8380,WX8381,
    WX8382,WX8383,WX8384,WX8385,WX8386,WX8387,WX8388,WX8389,WX8390,WX8391,
    WX8392,WX8393,WX8394,WX8395,WX8396,WX8397,WX8398,WX8399,WX8400,WX8401,
    WX8690,WX8674,WX8692,WX8675,WX8694,WX8676,WX8696,WX8677,WX8698,WX8678,
    WX8700,WX8679,WX8702,WX8680,WX8704,WX8681,WX8706,WX8682,WX8708,WX8683,
    WX8710,WX8684,WX8712,WX8685,WX8714,WX8686,WX8716,WX8687,WX8718,WX8688,
    WX8720,WX8689,WX8722,WX8658,WX8724,WX8659,WX8726,WX8660,WX8728,WX8661,
    WX8730,WX8662,WX8732,WX8663,WX8734,WX8664,WX8736,WX8665,WX8738,WX8666,
    WX8740,WX8667,WX8742,WX8668,WX8744,WX8669,WX8746,WX8670,WX8748,WX8671,
    WX8750,WX8672,WX8752,WX8673,WX8754,WX8755,WX8756,WX8757,WX8758,WX8759,
    WX8760,WX8763,WX8767,WX8769,WX8768,WX8770,WX8774,WX8776,WX8775,WX8777,
    WX8781,WX8783,WX8782,WX8784,WX8788,WX8790,WX8789,WX8791,WX8795,WX8797,
    WX8796,WX8798,WX8802,WX8804,WX8803,WX8805,WX8809,WX8811,WX8810,WX8812,
    WX8816,WX8818,WX8817,WX8819,WX8823,WX8825,WX8824,WX8826,WX8830,WX8832,
    WX8831,WX8833,WX8837,WX8839,WX8838,WX8840,WX8844,WX8846,WX8845,WX8847,
    WX8851,WX8853,WX8852,WX8854,WX8858,WX8860,WX8859,WX8861,WX8865,WX8867,
    WX8866,WX8868,WX8872,WX8874,WX8873,WX8875,WX8879,WX8881,WX8880,WX8882,
    WX8886,WX8888,WX8887,WX8889,WX8893,WX8895,WX8894,WX8896,WX8900,WX8902,
    WX8901,WX8903,WX8907,WX8909,WX8908,WX8910,WX8914,WX8916,WX8915,WX8917,
    WX8921,WX8923,WX8922,WX8924,WX8928,WX8930,WX8929,WX8931,WX8935,WX8937,
    WX8936,WX8938,WX8942,WX8944,WX8943,WX8945,WX8949,WX8951,WX8950,WX8952,
    WX8956,WX8958,WX8957,WX8959,WX8963,WX8965,WX8964,WX8966,WX8970,WX8972,
    WX8971,WX8973,WX8977,WX8979,WX8978,WX8980,WX8984,WX8986,WX8985,WX8987,
    WX8988,WX9021,WX9088,WX10054,WX9092,WX10055,WX9096,WX9098,WX9089,WX9099,
    WX9102,WX9106,WX9110,WX9112,WX9103,WX9113,WX9116,WX9120,WX9124,WX9126,
    WX9117,WX9127,WX9130,WX9134,WX9138,WX9140,WX9131,WX9141,WX9144,WX9148,
    WX9152,WX9154,WX9145,WX9155,WX9158,WX9162,WX9166,WX9168,WX9159,WX9169,
    WX9172,WX9176,WX9180,WX9182,WX9173,WX9183,WX9186,WX9190,WX9194,WX9196,
    WX9187,WX9197,WX9200,WX9204,WX9208,WX9210,WX9201,WX9211,WX9214,WX9218,
    WX9222,WX9224,WX9215,WX9225,WX9228,WX9232,WX9236,WX9238,WX9229,WX9239,
    WX9242,WX9246,WX9250,WX9252,WX9243,WX9253,WX9256,WX9260,WX9264,WX9266,
    WX9257,WX9267,WX9270,WX9274,WX9278,WX9280,WX9271,WX9281,WX9284,WX9288,
    WX9292,WX9294,WX9285,WX9295,WX9298,WX9302,WX9306,WX9308,WX9299,WX9309,
    WX9312,WX9316,WX9320,WX9322,WX9313,WX9323,WX9326,WX9330,WX9334,WX9336,
    WX9327,WX9337,WX9340,WX9344,WX9348,WX9350,WX9341,WX9351,WX9354,WX9358,
    WX9362,WX9364,WX9355,WX9365,WX9368,WX9372,WX9376,WX9378,WX9369,WX9379,
    WX9382,WX9386,WX9390,WX9392,WX9383,WX9393,WX9396,WX9400,WX9404,WX9406,
    WX9397,WX9407,WX9410,WX9414,WX9418,WX9420,WX9411,WX9421,WX9424,WX9428,
    WX9432,WX9434,WX9425,WX9435,WX9438,WX9442,WX9446,WX9448,WX9439,WX9449,
    WX9452,WX9456,WX9460,WX9462,WX9453,WX9463,WX9466,WX9470,WX9474,WX9476,
    WX9467,WX9477,WX9480,WX9484,WX9488,WX9490,WX9481,WX9491,WX9494,WX9498,
    WX9502,WX9504,WX9495,WX9505,WX9508,WX9512,WX9516,WX9518,WX9509,WX9519,
    WX9522,WX9526,WX9530,WX9532,WX9523,WX9533,WX9534,WX9599,WX10016,WX9600,
    WX10018,WX9601,WX10020,WX9602,WX10022,WX9603,WX10024,WX9604,WX10026,WX9605,
    WX10028,WX9606,WX10030,WX9607,WX10032,WX9608,WX10034,WX9609,WX10036,WX9610,
    WX10038,WX9611,WX10040,WX9612,WX10042,WX9613,WX10044,WX9614,WX10046,WX9615,
    WX9984,WX9616,WX9986,WX9617,WX9988,WX9618,WX9990,WX9619,WX9992,WX9620,
    WX9994,WX9621,WX9996,WX9622,WX9998,WX9623,WX10000,WX9624,WX10002,WX9625,
    WX10004,WX9626,WX10006,WX9627,WX10008,WX9628,WX10010,WX9629,WX10012,WX9630,
    WX10014,WX9631,WX9632,WX9633,WX9634,WX9635,WX9636,WX9637,WX9638,WX9639,
    WX9640,WX9641,WX9642,WX9643,WX9644,WX9645,WX9646,WX9647,WX9648,WX9649,
    WX9650,WX9651,WX9652,WX9653,WX9654,WX9655,WX9656,WX9657,WX9658,WX9659,
    WX9660,WX9661,WX9662,WX9663,WX9664,WX9665,WX9666,WX9667,WX9668,WX9669,
    WX9670,WX9671,WX9672,WX9673,WX9674,WX9675,WX9676,WX9677,WX9678,WX9679,
    WX9680,WX9681,WX9682,WX9683,WX9684,WX9685,WX9686,WX9687,WX9688,WX9689,
    WX9690,WX9691,WX9692,WX9693,WX9694,WX9983,WX9967,WX9985,WX9968,WX9987,
    WX9969,WX9989,WX9970,WX9991,WX9971,WX9993,WX9972,WX9995,WX9973,WX9997,
    WX9974,WX9999,WX9975,WX10001,WX9976,WX10003,WX9977,WX10005,WX9978,WX10007,
    WX9979,WX10009,WX9980,WX10011,WX9981,WX10013,WX9982,WX10015,WX9951,WX10017,
    WX9952,WX10019,WX9953,WX10021,WX9954,WX10023,WX9955,WX10025,WX9956,WX10027,
    WX9957,WX10029,WX9958,WX10031,WX9959,WX10033,WX9960,WX10035,WX9961,WX10037,
    WX9962,WX10039,WX9963,WX10041,WX9964,WX10043,WX9965,WX10045,WX9966,WX10047,
    WX10048,WX10049,WX10050,WX10051,WX10052,WX10053,WX10056,WX10060,WX10062,
    WX10061,WX10063,WX10067,WX10069,WX10068,WX10070,WX10074,WX10076,WX10075,
    WX10077,WX10081,WX10083,WX10082,WX10084,WX10088,WX10090,WX10089,WX10091,
    WX10095,WX10097,WX10096,WX10098,WX10102,WX10104,WX10103,WX10105,WX10109,
    WX10111,WX10110,WX10112,WX10116,WX10118,WX10117,WX10119,WX10123,WX10125,
    WX10124,WX10126,WX10130,WX10132,WX10131,WX10133,WX10137,WX10139,WX10138,
    WX10140,WX10144,WX10146,WX10145,WX10147,WX10151,WX10153,WX10152,WX10154,
    WX10158,WX10160,WX10159,WX10161,WX10165,WX10167,WX10166,WX10168,WX10172,
    WX10174,WX10173,WX10175,WX10179,WX10181,WX10180,WX10182,WX10186,WX10188,
    WX10187,WX10189,WX10193,WX10195,WX10194,WX10196,WX10200,WX10202,WX10201,
    WX10203,WX10207,WX10209,WX10208,WX10210,WX10214,WX10216,WX10215,WX10217,
    WX10221,WX10223,WX10222,WX10224,WX10228,WX10230,WX10229,WX10231,WX10235,
    WX10237,WX10236,WX10238,WX10242,WX10244,WX10243,WX10245,WX10249,WX10251,
    WX10250,WX10252,WX10256,WX10258,WX10257,WX10259,WX10263,WX10265,WX10264,
    WX10266,WX10270,WX10272,WX10271,WX10273,WX10277,WX10279,WX10278,WX10280,
    WX10281,WX10314,WX10381,WX11347,WX10385,WX11348,WX10389,WX10391,WX10382,
    WX10392,WX10395,WX10399,WX10403,WX10405,WX10396,WX10406,WX10409,WX10413,
    WX10417,WX10419,WX10410,WX10420,WX10423,WX10427,WX10431,WX10433,WX10424,
    WX10434,WX10437,WX10441,WX10445,WX10447,WX10438,WX10448,WX10451,WX10455,
    WX10459,WX10461,WX10452,WX10462,WX10465,WX10469,WX10473,WX10475,WX10466,
    WX10476,WX10479,WX10483,WX10487,WX10489,WX10480,WX10490,WX10493,WX10497,
    WX10501,WX10503,WX10494,WX10504,WX10507,WX10511,WX10515,WX10517,WX10508,
    WX10518,WX10521,WX10525,WX10529,WX10531,WX10522,WX10532,WX10535,WX10539,
    WX10543,WX10545,WX10536,WX10546,WX10549,WX10553,WX10557,WX10559,WX10550,
    WX10560,WX10563,WX10567,WX10571,WX10573,WX10564,WX10574,WX10577,WX10581,
    WX10585,WX10587,WX10578,WX10588,WX10591,WX10595,WX10599,WX10601,WX10592,
    WX10602,WX10605,WX10609,WX10613,WX10615,WX10606,WX10616,WX10619,WX10623,
    WX10627,WX10629,WX10620,WX10630,WX10633,WX10637,WX10641,WX10643,WX10634,
    WX10644,WX10647,WX10651,WX10655,WX10657,WX10648,WX10658,WX10661,WX10665,
    WX10669,WX10671,WX10662,WX10672,WX10675,WX10679,WX10683,WX10685,WX10676,
    WX10686,WX10689,WX10693,WX10697,WX10699,WX10690,WX10700,WX10703,WX10707,
    WX10711,WX10713,WX10704,WX10714,WX10717,WX10721,WX10725,WX10727,WX10718,
    WX10728,WX10731,WX10735,WX10739,WX10741,WX10732,WX10742,WX10745,WX10749,
    WX10753,WX10755,WX10746,WX10756,WX10759,WX10763,WX10767,WX10769,WX10760,
    WX10770,WX10773,WX10777,WX10781,WX10783,WX10774,WX10784,WX10787,WX10791,
    WX10795,WX10797,WX10788,WX10798,WX10801,WX10805,WX10809,WX10811,WX10802,
    WX10812,WX10815,WX10819,WX10823,WX10825,WX10816,WX10826,WX10827,WX10892,
    WX11309,WX10893,WX11311,WX10894,WX11313,WX10895,WX11315,WX10896,WX11317,
    WX10897,WX11319,WX10898,WX11321,WX10899,WX11323,WX10900,WX11325,WX10901,
    WX11327,WX10902,WX11329,WX10903,WX11331,WX10904,WX11333,WX10905,WX11335,
    WX10906,WX11337,WX10907,WX11339,WX10908,WX11277,WX10909,WX11279,WX10910,
    WX11281,WX10911,WX11283,WX10912,WX11285,WX10913,WX11287,WX10914,WX11289,
    WX10915,WX11291,WX10916,WX11293,WX10917,WX11295,WX10918,WX11297,WX10919,
    WX11299,WX10920,WX11301,WX10921,WX11303,WX10922,WX11305,WX10923,WX11307,
    WX10924,WX10925,WX10926,WX10927,WX10928,WX10929,WX10930,WX10931,WX10932,
    WX10933,WX10934,WX10935,WX10936,WX10937,WX10938,WX10939,WX10940,WX10941,
    WX10942,WX10943,WX10944,WX10945,WX10946,WX10947,WX10948,WX10949,WX10950,
    WX10951,WX10952,WX10953,WX10954,WX10955,WX10956,WX10957,WX10958,WX10959,
    WX10960,WX10961,WX10962,WX10963,WX10964,WX10965,WX10966,WX10967,WX10968,
    WX10969,WX10970,WX10971,WX10972,WX10973,WX10974,WX10975,WX10976,WX10977,
    WX10978,WX10979,WX10980,WX10981,WX10982,WX10983,WX10984,WX10985,WX10986,
    WX10987,WX11276,WX11260,WX11278,WX11261,WX11280,WX11262,WX11282,WX11263,
    WX11284,WX11264,WX11286,WX11265,WX11288,WX11266,WX11290,WX11267,WX11292,
    WX11268,WX11294,WX11269,WX11296,WX11270,WX11298,WX11271,WX11300,WX11272,
    WX11302,WX11273,WX11304,WX11274,WX11306,WX11275,WX11308,WX11244,WX11310,
    WX11245,WX11312,WX11246,WX11314,WX11247,WX11316,WX11248,WX11318,WX11249,
    WX11320,WX11250,WX11322,WX11251,WX11324,WX11252,WX11326,WX11253,WX11328,
    WX11254,WX11330,WX11255,WX11332,WX11256,WX11334,WX11257,WX11336,WX11258,
    WX11338,WX11259,WX11340,WX11341,WX11342,WX11343,WX11344,WX11345,WX11346,
    WX11349,WX11353,WX11355,WX11354,WX11356,WX11360,WX11362,WX11361,WX11363,
    WX11367,WX11369,WX11368,WX11370,WX11374,WX11376,WX11375,WX11377,WX11381,
    WX11383,WX11382,WX11384,WX11388,WX11390,WX11389,WX11391,WX11395,WX11397,
    WX11396,WX11398,WX11402,WX11404,WX11403,WX11405,WX11409,WX11411,WX11410,
    WX11412,WX11416,WX11418,WX11417,WX11419,WX11423,WX11425,WX11424,WX11426,
    WX11430,WX11432,WX11431,WX11433,WX11437,WX11439,WX11438,WX11440,WX11444,
    WX11446,WX11445,WX11447,WX11451,WX11453,WX11452,WX11454,WX11458,WX11460,
    WX11459,WX11461,WX11465,WX11467,WX11466,WX11468,WX11472,WX11474,WX11473,
    WX11475,WX11479,WX11481,WX11480,WX11482,WX11486,WX11488,WX11487,WX11489,
    WX11493,WX11495,WX11494,WX11496,WX11500,WX11502,WX11501,WX11503,WX11507,
    WX11509,WX11508,WX11510,WX11514,WX11516,WX11515,WX11517,WX11521,WX11523,
    WX11522,WX11524,WX11528,WX11530,WX11529,WX11531,WX11535,WX11537,WX11536,
    WX11538,WX11542,WX11544,WX11543,WX11545,WX11549,WX11551,WX11550,WX11552,
    WX11556,WX11558,WX11557,WX11559,WX11563,WX11565,WX11564,WX11566,WX11570,
    WX11572,WX11571,WX11573,WX11574,WX11607,WX35,WX46,WX36,WX42,WX39,WX40,WX43,
    WX44,WX49,WX60,WX50,WX56,WX53,WX54,WX57,WX58,WX63,WX74,WX64,WX70,WX67,WX68,
    WX71,WX72,WX77,WX88,WX78,WX84,WX81,WX82,WX85,WX86,WX91,WX102,WX92,WX98,
    WX95,WX96,WX99,WX100,WX105,WX116,WX106,WX112,WX109,WX110,WX113,WX114,WX119,
    WX130,WX120,WX126,WX123,WX124,WX127,WX128,WX133,WX144,WX134,WX140,WX137,
    WX138,WX141,WX142,WX147,WX158,WX148,WX154,WX151,WX152,WX155,WX156,WX161,
    WX172,WX162,WX168,WX165,WX166,WX169,WX170,WX175,WX186,WX176,WX182,WX179,
    WX180,WX183,WX184,WX189,WX200,WX190,WX196,WX193,WX194,WX197,WX198,WX203,
    WX214,WX204,WX210,WX207,WX208,WX211,WX212,WX217,WX228,WX218,WX224,WX221,
    WX222,WX225,WX226,WX231,WX242,WX232,WX238,WX235,WX236,WX239,WX240,WX245,
    WX256,WX246,WX252,WX249,WX250,WX253,WX254,WX259,WX270,WX260,WX266,WX263,
    WX264,WX267,WX268,WX273,WX284,WX274,WX280,WX277,WX278,WX281,WX282,WX287,
    WX298,WX288,WX294,WX291,WX292,WX295,WX296,WX301,WX312,WX302,WX308,WX305,
    WX306,WX309,WX310,WX315,WX326,WX316,WX322,WX319,WX320,WX323,WX324,WX329,
    WX340,WX330,WX336,WX333,WX334,WX337,WX338,WX343,WX354,WX344,WX350,WX347,
    WX348,WX351,WX352,WX357,WX368,WX358,WX364,WX361,WX362,WX365,WX366,WX371,
    WX382,WX372,WX378,WX375,WX376,WX379,WX380,WX385,WX396,WX386,WX392,WX389,
    WX390,WX393,WX394,WX399,WX410,WX400,WX406,WX403,WX404,WX407,WX408,WX413,
    WX424,WX414,WX420,WX417,WX418,WX421,WX422,WX427,WX438,WX428,WX434,WX431,
    WX432,WX435,WX436,WX441,WX452,WX442,WX448,WX445,WX446,WX449,WX450,WX455,
    WX466,WX456,WX462,WX459,WX460,WX463,WX464,WX469,WX480,WX470,WX476,WX473,
    WX474,WX477,WX478,WX1007,WX1006,WX1008,WX1014,WX1013,WX1015,WX1021,WX1020,
    WX1022,WX1028,WX1027,WX1029,WX1035,WX1034,WX1036,WX1042,WX1041,WX1043,
    WX1049,WX1048,WX1050,WX1056,WX1055,WX1057,WX1063,WX1062,WX1064,WX1070,
    WX1069,WX1071,WX1077,WX1076,WX1078,WX1084,WX1083,WX1085,WX1091,WX1090,
    WX1092,WX1098,WX1097,WX1099,WX1105,WX1104,WX1106,WX1112,WX1111,WX1113,
    WX1119,WX1118,WX1120,WX1126,WX1125,WX1127,WX1133,WX1132,WX1134,WX1140,
    WX1139,WX1141,WX1147,WX1146,WX1148,WX1154,WX1153,WX1155,WX1161,WX1160,
    WX1162,WX1168,WX1167,WX1169,WX1175,WX1174,WX1176,WX1182,WX1181,WX1183,
    WX1189,WX1188,WX1190,WX1196,WX1195,WX1197,WX1203,WX1202,WX1204,WX1210,
    WX1209,WX1211,WX1217,WX1216,WX1218,WX1224,WX1223,WX1225,WX1234,WX1262,
    WX1261,WX1260,WX1233,WX1259,WX1258,WX1257,WX1256,WX1255,WX1254,WX1232,
    WX1253,WX1252,WX1251,WX1250,WX1231,WX1249,WX1248,WX1247,WX1246,WX1245,
    WX1244,WX1243,WX1242,WX1241,WX1240,WX1239,WX1238,WX1237,WX1236,WX1235,
    WX1328,WX1339,WX1329,WX1335,WX1332,WX1333,WX1336,WX1337,WX1342,WX1353,
    WX1343,WX1349,WX1346,WX1347,WX1350,WX1351,WX1356,WX1367,WX1357,WX1363,
    WX1360,WX1361,WX1364,WX1365,WX1370,WX1381,WX1371,WX1377,WX1374,WX1375,
    WX1378,WX1379,WX1384,WX1395,WX1385,WX1391,WX1388,WX1389,WX1392,WX1393,
    WX1398,WX1409,WX1399,WX1405,WX1402,WX1403,WX1406,WX1407,WX1412,WX1423,
    WX1413,WX1419,WX1416,WX1417,WX1420,WX1421,WX1426,WX1437,WX1427,WX1433,
    WX1430,WX1431,WX1434,WX1435,WX1440,WX1451,WX1441,WX1447,WX1444,WX1445,
    WX1448,WX1449,WX1454,WX1465,WX1455,WX1461,WX1458,WX1459,WX1462,WX1463,
    WX1468,WX1479,WX1469,WX1475,WX1472,WX1473,WX1476,WX1477,WX1482,WX1493,
    WX1483,WX1489,WX1486,WX1487,WX1490,WX1491,WX1496,WX1507,WX1497,WX1503,
    WX1500,WX1501,WX1504,WX1505,WX1510,WX1521,WX1511,WX1517,WX1514,WX1515,
    WX1518,WX1519,WX1524,WX1535,WX1525,WX1531,WX1528,WX1529,WX1532,WX1533,
    WX1538,WX1549,WX1539,WX1545,WX1542,WX1543,WX1546,WX1547,WX1552,WX1563,
    WX1553,WX1559,WX1556,WX1557,WX1560,WX1561,WX1566,WX1577,WX1567,WX1573,
    WX1570,WX1571,WX1574,WX1575,WX1580,WX1591,WX1581,WX1587,WX1584,WX1585,
    WX1588,WX1589,WX1594,WX1605,WX1595,WX1601,WX1598,WX1599,WX1602,WX1603,
    WX1608,WX1619,WX1609,WX1615,WX1612,WX1613,WX1616,WX1617,WX1622,WX1633,
    WX1623,WX1629,WX1626,WX1627,WX1630,WX1631,WX1636,WX1647,WX1637,WX1643,
    WX1640,WX1641,WX1644,WX1645,WX1650,WX1661,WX1651,WX1657,WX1654,WX1655,
    WX1658,WX1659,WX1664,WX1675,WX1665,WX1671,WX1668,WX1669,WX1672,WX1673,
    WX1678,WX1689,WX1679,WX1685,WX1682,WX1683,WX1686,WX1687,WX1692,WX1703,
    WX1693,WX1699,WX1696,WX1697,WX1700,WX1701,WX1706,WX1717,WX1707,WX1713,
    WX1710,WX1711,WX1714,WX1715,WX1720,WX1731,WX1721,WX1727,WX1724,WX1725,
    WX1728,WX1729,WX1734,WX1745,WX1735,WX1741,WX1738,WX1739,WX1742,WX1743,
    WX1748,WX1759,WX1749,WX1755,WX1752,WX1753,WX1756,WX1757,WX1762,WX1773,
    WX1763,WX1769,WX1766,WX1767,WX1770,WX1771,WX2300,WX2299,WX2301,WX2307,
    WX2306,WX2308,WX2314,WX2313,WX2315,WX2321,WX2320,WX2322,WX2328,WX2327,
    WX2329,WX2335,WX2334,WX2336,WX2342,WX2341,WX2343,WX2349,WX2348,WX2350,
    WX2356,WX2355,WX2357,WX2363,WX2362,WX2364,WX2370,WX2369,WX2371,WX2377,
    WX2376,WX2378,WX2384,WX2383,WX2385,WX2391,WX2390,WX2392,WX2398,WX2397,
    WX2399,WX2405,WX2404,WX2406,WX2412,WX2411,WX2413,WX2419,WX2418,WX2420,
    WX2426,WX2425,WX2427,WX2433,WX2432,WX2434,WX2440,WX2439,WX2441,WX2447,
    WX2446,WX2448,WX2454,WX2453,WX2455,WX2461,WX2460,WX2462,WX2468,WX2467,
    WX2469,WX2475,WX2474,WX2476,WX2482,WX2481,WX2483,WX2489,WX2488,WX2490,
    WX2496,WX2495,WX2497,WX2503,WX2502,WX2504,WX2510,WX2509,WX2511,WX2517,
    WX2516,WX2518,WX2527,WX2555,WX2554,WX2553,WX2526,WX2552,WX2551,WX2550,
    WX2549,WX2548,WX2547,WX2525,WX2546,WX2545,WX2544,WX2543,WX2524,WX2542,
    WX2541,WX2540,WX2539,WX2538,WX2537,WX2536,WX2535,WX2534,WX2533,WX2532,
    WX2531,WX2530,WX2529,WX2528,WX2621,WX2632,WX2622,WX2628,WX2625,WX2626,
    WX2629,WX2630,WX2635,WX2646,WX2636,WX2642,WX2639,WX2640,WX2643,WX2644,
    WX2649,WX2660,WX2650,WX2656,WX2653,WX2654,WX2657,WX2658,WX2663,WX2674,
    WX2664,WX2670,WX2667,WX2668,WX2671,WX2672,WX2677,WX2688,WX2678,WX2684,
    WX2681,WX2682,WX2685,WX2686,WX2691,WX2702,WX2692,WX2698,WX2695,WX2696,
    WX2699,WX2700,WX2705,WX2716,WX2706,WX2712,WX2709,WX2710,WX2713,WX2714,
    WX2719,WX2730,WX2720,WX2726,WX2723,WX2724,WX2727,WX2728,WX2733,WX2744,
    WX2734,WX2740,WX2737,WX2738,WX2741,WX2742,WX2747,WX2758,WX2748,WX2754,
    WX2751,WX2752,WX2755,WX2756,WX2761,WX2772,WX2762,WX2768,WX2765,WX2766,
    WX2769,WX2770,WX2775,WX2786,WX2776,WX2782,WX2779,WX2780,WX2783,WX2784,
    WX2789,WX2800,WX2790,WX2796,WX2793,WX2794,WX2797,WX2798,WX2803,WX2814,
    WX2804,WX2810,WX2807,WX2808,WX2811,WX2812,WX2817,WX2828,WX2818,WX2824,
    WX2821,WX2822,WX2825,WX2826,WX2831,WX2842,WX2832,WX2838,WX2835,WX2836,
    WX2839,WX2840,WX2845,WX2856,WX2846,WX2852,WX2849,WX2850,WX2853,WX2854,
    WX2859,WX2870,WX2860,WX2866,WX2863,WX2864,WX2867,WX2868,WX2873,WX2884,
    WX2874,WX2880,WX2877,WX2878,WX2881,WX2882,WX2887,WX2898,WX2888,WX2894,
    WX2891,WX2892,WX2895,WX2896,WX2901,WX2912,WX2902,WX2908,WX2905,WX2906,
    WX2909,WX2910,WX2915,WX2926,WX2916,WX2922,WX2919,WX2920,WX2923,WX2924,
    WX2929,WX2940,WX2930,WX2936,WX2933,WX2934,WX2937,WX2938,WX2943,WX2954,
    WX2944,WX2950,WX2947,WX2948,WX2951,WX2952,WX2957,WX2968,WX2958,WX2964,
    WX2961,WX2962,WX2965,WX2966,WX2971,WX2982,WX2972,WX2978,WX2975,WX2976,
    WX2979,WX2980,WX2985,WX2996,WX2986,WX2992,WX2989,WX2990,WX2993,WX2994,
    WX2999,WX3010,WX3000,WX3006,WX3003,WX3004,WX3007,WX3008,WX3013,WX3024,
    WX3014,WX3020,WX3017,WX3018,WX3021,WX3022,WX3027,WX3038,WX3028,WX3034,
    WX3031,WX3032,WX3035,WX3036,WX3041,WX3052,WX3042,WX3048,WX3045,WX3046,
    WX3049,WX3050,WX3055,WX3066,WX3056,WX3062,WX3059,WX3060,WX3063,WX3064,
    WX3593,WX3592,WX3594,WX3600,WX3599,WX3601,WX3607,WX3606,WX3608,WX3614,
    WX3613,WX3615,WX3621,WX3620,WX3622,WX3628,WX3627,WX3629,WX3635,WX3634,
    WX3636,WX3642,WX3641,WX3643,WX3649,WX3648,WX3650,WX3656,WX3655,WX3657,
    WX3663,WX3662,WX3664,WX3670,WX3669,WX3671,WX3677,WX3676,WX3678,WX3684,
    WX3683,WX3685,WX3691,WX3690,WX3692,WX3698,WX3697,WX3699,WX3705,WX3704,
    WX3706,WX3712,WX3711,WX3713,WX3719,WX3718,WX3720,WX3726,WX3725,WX3727,
    WX3733,WX3732,WX3734,WX3740,WX3739,WX3741,WX3747,WX3746,WX3748,WX3754,
    WX3753,WX3755,WX3761,WX3760,WX3762,WX3768,WX3767,WX3769,WX3775,WX3774,
    WX3776,WX3782,WX3781,WX3783,WX3789,WX3788,WX3790,WX3796,WX3795,WX3797,
    WX3803,WX3802,WX3804,WX3810,WX3809,WX3811,WX3820,WX3848,WX3847,WX3846,
    WX3819,WX3845,WX3844,WX3843,WX3842,WX3841,WX3840,WX3818,WX3839,WX3838,
    WX3837,WX3836,WX3817,WX3835,WX3834,WX3833,WX3832,WX3831,WX3830,WX3829,
    WX3828,WX3827,WX3826,WX3825,WX3824,WX3823,WX3822,WX3821,WX3914,WX3925,
    WX3915,WX3921,WX3918,WX3919,WX3922,WX3923,WX3928,WX3939,WX3929,WX3935,
    WX3932,WX3933,WX3936,WX3937,WX3942,WX3953,WX3943,WX3949,WX3946,WX3947,
    WX3950,WX3951,WX3956,WX3967,WX3957,WX3963,WX3960,WX3961,WX3964,WX3965,
    WX3970,WX3981,WX3971,WX3977,WX3974,WX3975,WX3978,WX3979,WX3984,WX3995,
    WX3985,WX3991,WX3988,WX3989,WX3992,WX3993,WX3998,WX4009,WX3999,WX4005,
    WX4002,WX4003,WX4006,WX4007,WX4012,WX4023,WX4013,WX4019,WX4016,WX4017,
    WX4020,WX4021,WX4026,WX4037,WX4027,WX4033,WX4030,WX4031,WX4034,WX4035,
    WX4040,WX4051,WX4041,WX4047,WX4044,WX4045,WX4048,WX4049,WX4054,WX4065,
    WX4055,WX4061,WX4058,WX4059,WX4062,WX4063,WX4068,WX4079,WX4069,WX4075,
    WX4072,WX4073,WX4076,WX4077,WX4082,WX4093,WX4083,WX4089,WX4086,WX4087,
    WX4090,WX4091,WX4096,WX4107,WX4097,WX4103,WX4100,WX4101,WX4104,WX4105,
    WX4110,WX4121,WX4111,WX4117,WX4114,WX4115,WX4118,WX4119,WX4124,WX4135,
    WX4125,WX4131,WX4128,WX4129,WX4132,WX4133,WX4138,WX4149,WX4139,WX4145,
    WX4142,WX4143,WX4146,WX4147,WX4152,WX4163,WX4153,WX4159,WX4156,WX4157,
    WX4160,WX4161,WX4166,WX4177,WX4167,WX4173,WX4170,WX4171,WX4174,WX4175,
    WX4180,WX4191,WX4181,WX4187,WX4184,WX4185,WX4188,WX4189,WX4194,WX4205,
    WX4195,WX4201,WX4198,WX4199,WX4202,WX4203,WX4208,WX4219,WX4209,WX4215,
    WX4212,WX4213,WX4216,WX4217,WX4222,WX4233,WX4223,WX4229,WX4226,WX4227,
    WX4230,WX4231,WX4236,WX4247,WX4237,WX4243,WX4240,WX4241,WX4244,WX4245,
    WX4250,WX4261,WX4251,WX4257,WX4254,WX4255,WX4258,WX4259,WX4264,WX4275,
    WX4265,WX4271,WX4268,WX4269,WX4272,WX4273,WX4278,WX4289,WX4279,WX4285,
    WX4282,WX4283,WX4286,WX4287,WX4292,WX4303,WX4293,WX4299,WX4296,WX4297,
    WX4300,WX4301,WX4306,WX4317,WX4307,WX4313,WX4310,WX4311,WX4314,WX4315,
    WX4320,WX4331,WX4321,WX4327,WX4324,WX4325,WX4328,WX4329,WX4334,WX4345,
    WX4335,WX4341,WX4338,WX4339,WX4342,WX4343,WX4348,WX4359,WX4349,WX4355,
    WX4352,WX4353,WX4356,WX4357,WX4886,WX4885,WX4887,WX4893,WX4892,WX4894,
    WX4900,WX4899,WX4901,WX4907,WX4906,WX4908,WX4914,WX4913,WX4915,WX4921,
    WX4920,WX4922,WX4928,WX4927,WX4929,WX4935,WX4934,WX4936,WX4942,WX4941,
    WX4943,WX4949,WX4948,WX4950,WX4956,WX4955,WX4957,WX4963,WX4962,WX4964,
    WX4970,WX4969,WX4971,WX4977,WX4976,WX4978,WX4984,WX4983,WX4985,WX4991,
    WX4990,WX4992,WX4998,WX4997,WX4999,WX5005,WX5004,WX5006,WX5012,WX5011,
    WX5013,WX5019,WX5018,WX5020,WX5026,WX5025,WX5027,WX5033,WX5032,WX5034,
    WX5040,WX5039,WX5041,WX5047,WX5046,WX5048,WX5054,WX5053,WX5055,WX5061,
    WX5060,WX5062,WX5068,WX5067,WX5069,WX5075,WX5074,WX5076,WX5082,WX5081,
    WX5083,WX5089,WX5088,WX5090,WX5096,WX5095,WX5097,WX5103,WX5102,WX5104,
    WX5113,WX5141,WX5140,WX5139,WX5112,WX5138,WX5137,WX5136,WX5135,WX5134,
    WX5133,WX5111,WX5132,WX5131,WX5130,WX5129,WX5110,WX5128,WX5127,WX5126,
    WX5125,WX5124,WX5123,WX5122,WX5121,WX5120,WX5119,WX5118,WX5117,WX5116,
    WX5115,WX5114,WX5207,WX5218,WX5208,WX5214,WX5211,WX5212,WX5215,WX5216,
    WX5221,WX5232,WX5222,WX5228,WX5225,WX5226,WX5229,WX5230,WX5235,WX5246,
    WX5236,WX5242,WX5239,WX5240,WX5243,WX5244,WX5249,WX5260,WX5250,WX5256,
    WX5253,WX5254,WX5257,WX5258,WX5263,WX5274,WX5264,WX5270,WX5267,WX5268,
    WX5271,WX5272,WX5277,WX5288,WX5278,WX5284,WX5281,WX5282,WX5285,WX5286,
    WX5291,WX5302,WX5292,WX5298,WX5295,WX5296,WX5299,WX5300,WX5305,WX5316,
    WX5306,WX5312,WX5309,WX5310,WX5313,WX5314,WX5319,WX5330,WX5320,WX5326,
    WX5323,WX5324,WX5327,WX5328,WX5333,WX5344,WX5334,WX5340,WX5337,WX5338,
    WX5341,WX5342,WX5347,WX5358,WX5348,WX5354,WX5351,WX5352,WX5355,WX5356,
    WX5361,WX5372,WX5362,WX5368,WX5365,WX5366,WX5369,WX5370,WX5375,WX5386,
    WX5376,WX5382,WX5379,WX5380,WX5383,WX5384,WX5389,WX5400,WX5390,WX5396,
    WX5393,WX5394,WX5397,WX5398,WX5403,WX5414,WX5404,WX5410,WX5407,WX5408,
    WX5411,WX5412,WX5417,WX5428,WX5418,WX5424,WX5421,WX5422,WX5425,WX5426,
    WX5431,WX5442,WX5432,WX5438,WX5435,WX5436,WX5439,WX5440,WX5445,WX5456,
    WX5446,WX5452,WX5449,WX5450,WX5453,WX5454,WX5459,WX5470,WX5460,WX5466,
    WX5463,WX5464,WX5467,WX5468,WX5473,WX5484,WX5474,WX5480,WX5477,WX5478,
    WX5481,WX5482,WX5487,WX5498,WX5488,WX5494,WX5491,WX5492,WX5495,WX5496,
    WX5501,WX5512,WX5502,WX5508,WX5505,WX5506,WX5509,WX5510,WX5515,WX5526,
    WX5516,WX5522,WX5519,WX5520,WX5523,WX5524,WX5529,WX5540,WX5530,WX5536,
    WX5533,WX5534,WX5537,WX5538,WX5543,WX5554,WX5544,WX5550,WX5547,WX5548,
    WX5551,WX5552,WX5557,WX5568,WX5558,WX5564,WX5561,WX5562,WX5565,WX5566,
    WX5571,WX5582,WX5572,WX5578,WX5575,WX5576,WX5579,WX5580,WX5585,WX5596,
    WX5586,WX5592,WX5589,WX5590,WX5593,WX5594,WX5599,WX5610,WX5600,WX5606,
    WX5603,WX5604,WX5607,WX5608,WX5613,WX5624,WX5614,WX5620,WX5617,WX5618,
    WX5621,WX5622,WX5627,WX5638,WX5628,WX5634,WX5631,WX5632,WX5635,WX5636,
    WX5641,WX5652,WX5642,WX5648,WX5645,WX5646,WX5649,WX5650,WX6179,WX6178,
    WX6180,WX6186,WX6185,WX6187,WX6193,WX6192,WX6194,WX6200,WX6199,WX6201,
    WX6207,WX6206,WX6208,WX6214,WX6213,WX6215,WX6221,WX6220,WX6222,WX6228,
    WX6227,WX6229,WX6235,WX6234,WX6236,WX6242,WX6241,WX6243,WX6249,WX6248,
    WX6250,WX6256,WX6255,WX6257,WX6263,WX6262,WX6264,WX6270,WX6269,WX6271,
    WX6277,WX6276,WX6278,WX6284,WX6283,WX6285,WX6291,WX6290,WX6292,WX6298,
    WX6297,WX6299,WX6305,WX6304,WX6306,WX6312,WX6311,WX6313,WX6319,WX6318,
    WX6320,WX6326,WX6325,WX6327,WX6333,WX6332,WX6334,WX6340,WX6339,WX6341,
    WX6347,WX6346,WX6348,WX6354,WX6353,WX6355,WX6361,WX6360,WX6362,WX6368,
    WX6367,WX6369,WX6375,WX6374,WX6376,WX6382,WX6381,WX6383,WX6389,WX6388,
    WX6390,WX6396,WX6395,WX6397,WX6406,WX6434,WX6433,WX6432,WX6405,WX6431,
    WX6430,WX6429,WX6428,WX6427,WX6426,WX6404,WX6425,WX6424,WX6423,WX6422,
    WX6403,WX6421,WX6420,WX6419,WX6418,WX6417,WX6416,WX6415,WX6414,WX6413,
    WX6412,WX6411,WX6410,WX6409,WX6408,WX6407,WX6500,WX6511,WX6501,WX6507,
    WX6504,WX6505,WX6508,WX6509,WX6514,WX6525,WX6515,WX6521,WX6518,WX6519,
    WX6522,WX6523,WX6528,WX6539,WX6529,WX6535,WX6532,WX6533,WX6536,WX6537,
    WX6542,WX6553,WX6543,WX6549,WX6546,WX6547,WX6550,WX6551,WX6556,WX6567,
    WX6557,WX6563,WX6560,WX6561,WX6564,WX6565,WX6570,WX6581,WX6571,WX6577,
    WX6574,WX6575,WX6578,WX6579,WX6584,WX6595,WX6585,WX6591,WX6588,WX6589,
    WX6592,WX6593,WX6598,WX6609,WX6599,WX6605,WX6602,WX6603,WX6606,WX6607,
    WX6612,WX6623,WX6613,WX6619,WX6616,WX6617,WX6620,WX6621,WX6626,WX6637,
    WX6627,WX6633,WX6630,WX6631,WX6634,WX6635,WX6640,WX6651,WX6641,WX6647,
    WX6644,WX6645,WX6648,WX6649,WX6654,WX6665,WX6655,WX6661,WX6658,WX6659,
    WX6662,WX6663,WX6668,WX6679,WX6669,WX6675,WX6672,WX6673,WX6676,WX6677,
    WX6682,WX6693,WX6683,WX6689,WX6686,WX6687,WX6690,WX6691,WX6696,WX6707,
    WX6697,WX6703,WX6700,WX6701,WX6704,WX6705,WX6710,WX6721,WX6711,WX6717,
    WX6714,WX6715,WX6718,WX6719,WX6724,WX6735,WX6725,WX6731,WX6728,WX6729,
    WX6732,WX6733,WX6738,WX6749,WX6739,WX6745,WX6742,WX6743,WX6746,WX6747,
    WX6752,WX6763,WX6753,WX6759,WX6756,WX6757,WX6760,WX6761,WX6766,WX6777,
    WX6767,WX6773,WX6770,WX6771,WX6774,WX6775,WX6780,WX6791,WX6781,WX6787,
    WX6784,WX6785,WX6788,WX6789,WX6794,WX6805,WX6795,WX6801,WX6798,WX6799,
    WX6802,WX6803,WX6808,WX6819,WX6809,WX6815,WX6812,WX6813,WX6816,WX6817,
    WX6822,WX6833,WX6823,WX6829,WX6826,WX6827,WX6830,WX6831,WX6836,WX6847,
    WX6837,WX6843,WX6840,WX6841,WX6844,WX6845,WX6850,WX6861,WX6851,WX6857,
    WX6854,WX6855,WX6858,WX6859,WX6864,WX6875,WX6865,WX6871,WX6868,WX6869,
    WX6872,WX6873,WX6878,WX6889,WX6879,WX6885,WX6882,WX6883,WX6886,WX6887,
    WX6892,WX6903,WX6893,WX6899,WX6896,WX6897,WX6900,WX6901,WX6906,WX6917,
    WX6907,WX6913,WX6910,WX6911,WX6914,WX6915,WX6920,WX6931,WX6921,WX6927,
    WX6924,WX6925,WX6928,WX6929,WX6934,WX6945,WX6935,WX6941,WX6938,WX6939,
    WX6942,WX6943,WX7472,WX7471,WX7473,WX7479,WX7478,WX7480,WX7486,WX7485,
    WX7487,WX7493,WX7492,WX7494,WX7500,WX7499,WX7501,WX7507,WX7506,WX7508,
    WX7514,WX7513,WX7515,WX7521,WX7520,WX7522,WX7528,WX7527,WX7529,WX7535,
    WX7534,WX7536,WX7542,WX7541,WX7543,WX7549,WX7548,WX7550,WX7556,WX7555,
    WX7557,WX7563,WX7562,WX7564,WX7570,WX7569,WX7571,WX7577,WX7576,WX7578,
    WX7584,WX7583,WX7585,WX7591,WX7590,WX7592,WX7598,WX7597,WX7599,WX7605,
    WX7604,WX7606,WX7612,WX7611,WX7613,WX7619,WX7618,WX7620,WX7626,WX7625,
    WX7627,WX7633,WX7632,WX7634,WX7640,WX7639,WX7641,WX7647,WX7646,WX7648,
    WX7654,WX7653,WX7655,WX7661,WX7660,WX7662,WX7668,WX7667,WX7669,WX7675,
    WX7674,WX7676,WX7682,WX7681,WX7683,WX7689,WX7688,WX7690,WX7699,WX7727,
    WX7726,WX7725,WX7698,WX7724,WX7723,WX7722,WX7721,WX7720,WX7719,WX7697,
    WX7718,WX7717,WX7716,WX7715,WX7696,WX7714,WX7713,WX7712,WX7711,WX7710,
    WX7709,WX7708,WX7707,WX7706,WX7705,WX7704,WX7703,WX7702,WX7701,WX7700,
    WX7793,WX7804,WX7794,WX7800,WX7797,WX7798,WX7801,WX7802,WX7807,WX7818,
    WX7808,WX7814,WX7811,WX7812,WX7815,WX7816,WX7821,WX7832,WX7822,WX7828,
    WX7825,WX7826,WX7829,WX7830,WX7835,WX7846,WX7836,WX7842,WX7839,WX7840,
    WX7843,WX7844,WX7849,WX7860,WX7850,WX7856,WX7853,WX7854,WX7857,WX7858,
    WX7863,WX7874,WX7864,WX7870,WX7867,WX7868,WX7871,WX7872,WX7877,WX7888,
    WX7878,WX7884,WX7881,WX7882,WX7885,WX7886,WX7891,WX7902,WX7892,WX7898,
    WX7895,WX7896,WX7899,WX7900,WX7905,WX7916,WX7906,WX7912,WX7909,WX7910,
    WX7913,WX7914,WX7919,WX7930,WX7920,WX7926,WX7923,WX7924,WX7927,WX7928,
    WX7933,WX7944,WX7934,WX7940,WX7937,WX7938,WX7941,WX7942,WX7947,WX7958,
    WX7948,WX7954,WX7951,WX7952,WX7955,WX7956,WX7961,WX7972,WX7962,WX7968,
    WX7965,WX7966,WX7969,WX7970,WX7975,WX7986,WX7976,WX7982,WX7979,WX7980,
    WX7983,WX7984,WX7989,WX8000,WX7990,WX7996,WX7993,WX7994,WX7997,WX7998,
    WX8003,WX8014,WX8004,WX8010,WX8007,WX8008,WX8011,WX8012,WX8017,WX8028,
    WX8018,WX8024,WX8021,WX8022,WX8025,WX8026,WX8031,WX8042,WX8032,WX8038,
    WX8035,WX8036,WX8039,WX8040,WX8045,WX8056,WX8046,WX8052,WX8049,WX8050,
    WX8053,WX8054,WX8059,WX8070,WX8060,WX8066,WX8063,WX8064,WX8067,WX8068,
    WX8073,WX8084,WX8074,WX8080,WX8077,WX8078,WX8081,WX8082,WX8087,WX8098,
    WX8088,WX8094,WX8091,WX8092,WX8095,WX8096,WX8101,WX8112,WX8102,WX8108,
    WX8105,WX8106,WX8109,WX8110,WX8115,WX8126,WX8116,WX8122,WX8119,WX8120,
    WX8123,WX8124,WX8129,WX8140,WX8130,WX8136,WX8133,WX8134,WX8137,WX8138,
    WX8143,WX8154,WX8144,WX8150,WX8147,WX8148,WX8151,WX8152,WX8157,WX8168,
    WX8158,WX8164,WX8161,WX8162,WX8165,WX8166,WX8171,WX8182,WX8172,WX8178,
    WX8175,WX8176,WX8179,WX8180,WX8185,WX8196,WX8186,WX8192,WX8189,WX8190,
    WX8193,WX8194,WX8199,WX8210,WX8200,WX8206,WX8203,WX8204,WX8207,WX8208,
    WX8213,WX8224,WX8214,WX8220,WX8217,WX8218,WX8221,WX8222,WX8227,WX8238,
    WX8228,WX8234,WX8231,WX8232,WX8235,WX8236,WX8765,WX8764,WX8766,WX8772,
    WX8771,WX8773,WX8779,WX8778,WX8780,WX8786,WX8785,WX8787,WX8793,WX8792,
    WX8794,WX8800,WX8799,WX8801,WX8807,WX8806,WX8808,WX8814,WX8813,WX8815,
    WX8821,WX8820,WX8822,WX8828,WX8827,WX8829,WX8835,WX8834,WX8836,WX8842,
    WX8841,WX8843,WX8849,WX8848,WX8850,WX8856,WX8855,WX8857,WX8863,WX8862,
    WX8864,WX8870,WX8869,WX8871,WX8877,WX8876,WX8878,WX8884,WX8883,WX8885,
    WX8891,WX8890,WX8892,WX8898,WX8897,WX8899,WX8905,WX8904,WX8906,WX8912,
    WX8911,WX8913,WX8919,WX8918,WX8920,WX8926,WX8925,WX8927,WX8933,WX8932,
    WX8934,WX8940,WX8939,WX8941,WX8947,WX8946,WX8948,WX8954,WX8953,WX8955,
    WX8961,WX8960,WX8962,WX8968,WX8967,WX8969,WX8975,WX8974,WX8976,WX8982,
    WX8981,WX8983,WX8992,WX9020,WX9019,WX9018,WX8991,WX9017,WX9016,WX9015,
    WX9014,WX9013,WX9012,WX8990,WX9011,WX9010,WX9009,WX9008,WX8989,WX9007,
    WX9006,WX9005,WX9004,WX9003,WX9002,WX9001,WX9000,WX8999,WX8998,WX8997,
    WX8996,WX8995,WX8994,WX8993,WX9086,WX9097,WX9087,WX9093,WX9090,WX9091,
    WX9094,WX9095,WX9100,WX9111,WX9101,WX9107,WX9104,WX9105,WX9108,WX9109,
    WX9114,WX9125,WX9115,WX9121,WX9118,WX9119,WX9122,WX9123,WX9128,WX9139,
    WX9129,WX9135,WX9132,WX9133,WX9136,WX9137,WX9142,WX9153,WX9143,WX9149,
    WX9146,WX9147,WX9150,WX9151,WX9156,WX9167,WX9157,WX9163,WX9160,WX9161,
    WX9164,WX9165,WX9170,WX9181,WX9171,WX9177,WX9174,WX9175,WX9178,WX9179,
    WX9184,WX9195,WX9185,WX9191,WX9188,WX9189,WX9192,WX9193,WX9198,WX9209,
    WX9199,WX9205,WX9202,WX9203,WX9206,WX9207,WX9212,WX9223,WX9213,WX9219,
    WX9216,WX9217,WX9220,WX9221,WX9226,WX9237,WX9227,WX9233,WX9230,WX9231,
    WX9234,WX9235,WX9240,WX9251,WX9241,WX9247,WX9244,WX9245,WX9248,WX9249,
    WX9254,WX9265,WX9255,WX9261,WX9258,WX9259,WX9262,WX9263,WX9268,WX9279,
    WX9269,WX9275,WX9272,WX9273,WX9276,WX9277,WX9282,WX9293,WX9283,WX9289,
    WX9286,WX9287,WX9290,WX9291,WX9296,WX9307,WX9297,WX9303,WX9300,WX9301,
    WX9304,WX9305,WX9310,WX9321,WX9311,WX9317,WX9314,WX9315,WX9318,WX9319,
    WX9324,WX9335,WX9325,WX9331,WX9328,WX9329,WX9332,WX9333,WX9338,WX9349,
    WX9339,WX9345,WX9342,WX9343,WX9346,WX9347,WX9352,WX9363,WX9353,WX9359,
    WX9356,WX9357,WX9360,WX9361,WX9366,WX9377,WX9367,WX9373,WX9370,WX9371,
    WX9374,WX9375,WX9380,WX9391,WX9381,WX9387,WX9384,WX9385,WX9388,WX9389,
    WX9394,WX9405,WX9395,WX9401,WX9398,WX9399,WX9402,WX9403,WX9408,WX9419,
    WX9409,WX9415,WX9412,WX9413,WX9416,WX9417,WX9422,WX9433,WX9423,WX9429,
    WX9426,WX9427,WX9430,WX9431,WX9436,WX9447,WX9437,WX9443,WX9440,WX9441,
    WX9444,WX9445,WX9450,WX9461,WX9451,WX9457,WX9454,WX9455,WX9458,WX9459,
    WX9464,WX9475,WX9465,WX9471,WX9468,WX9469,WX9472,WX9473,WX9478,WX9489,
    WX9479,WX9485,WX9482,WX9483,WX9486,WX9487,WX9492,WX9503,WX9493,WX9499,
    WX9496,WX9497,WX9500,WX9501,WX9506,WX9517,WX9507,WX9513,WX9510,WX9511,
    WX9514,WX9515,WX9520,WX9531,WX9521,WX9527,WX9524,WX9525,WX9528,WX9529,
    WX10058,WX10057,WX10059,WX10065,WX10064,WX10066,WX10072,WX10071,WX10073,
    WX10079,WX10078,WX10080,WX10086,WX10085,WX10087,WX10093,WX10092,WX10094,
    WX10100,WX10099,WX10101,WX10107,WX10106,WX10108,WX10114,WX10113,WX10115,
    WX10121,WX10120,WX10122,WX10128,WX10127,WX10129,WX10135,WX10134,WX10136,
    WX10142,WX10141,WX10143,WX10149,WX10148,WX10150,WX10156,WX10155,WX10157,
    WX10163,WX10162,WX10164,WX10170,WX10169,WX10171,WX10177,WX10176,WX10178,
    WX10184,WX10183,WX10185,WX10191,WX10190,WX10192,WX10198,WX10197,WX10199,
    WX10205,WX10204,WX10206,WX10212,WX10211,WX10213,WX10219,WX10218,WX10220,
    WX10226,WX10225,WX10227,WX10233,WX10232,WX10234,WX10240,WX10239,WX10241,
    WX10247,WX10246,WX10248,WX10254,WX10253,WX10255,WX10261,WX10260,WX10262,
    WX10268,WX10267,WX10269,WX10275,WX10274,WX10276,WX10285,WX10313,WX10312,
    WX10311,WX10284,WX10310,WX10309,WX10308,WX10307,WX10306,WX10305,WX10283,
    WX10304,WX10303,WX10302,WX10301,WX10282,WX10300,WX10299,WX10298,WX10297,
    WX10296,WX10295,WX10294,WX10293,WX10292,WX10291,WX10290,WX10289,WX10288,
    WX10287,WX10286,WX10379,WX10390,WX10380,WX10386,WX10383,WX10384,WX10387,
    WX10388,WX10393,WX10404,WX10394,WX10400,WX10397,WX10398,WX10401,WX10402,
    WX10407,WX10418,WX10408,WX10414,WX10411,WX10412,WX10415,WX10416,WX10421,
    WX10432,WX10422,WX10428,WX10425,WX10426,WX10429,WX10430,WX10435,WX10446,
    WX10436,WX10442,WX10439,WX10440,WX10443,WX10444,WX10449,WX10460,WX10450,
    WX10456,WX10453,WX10454,WX10457,WX10458,WX10463,WX10474,WX10464,WX10470,
    WX10467,WX10468,WX10471,WX10472,WX10477,WX10488,WX10478,WX10484,WX10481,
    WX10482,WX10485,WX10486,WX10491,WX10502,WX10492,WX10498,WX10495,WX10496,
    WX10499,WX10500,WX10505,WX10516,WX10506,WX10512,WX10509,WX10510,WX10513,
    WX10514,WX10519,WX10530,WX10520,WX10526,WX10523,WX10524,WX10527,WX10528,
    WX10533,WX10544,WX10534,WX10540,WX10537,WX10538,WX10541,WX10542,WX10547,
    WX10558,WX10548,WX10554,WX10551,WX10552,WX10555,WX10556,WX10561,WX10572,
    WX10562,WX10568,WX10565,WX10566,WX10569,WX10570,WX10575,WX10586,WX10576,
    WX10582,WX10579,WX10580,WX10583,WX10584,WX10589,WX10600,WX10590,WX10596,
    WX10593,WX10594,WX10597,WX10598,WX10603,WX10614,WX10604,WX10610,WX10607,
    WX10608,WX10611,WX10612,WX10617,WX10628,WX10618,WX10624,WX10621,WX10622,
    WX10625,WX10626,WX10631,WX10642,WX10632,WX10638,WX10635,WX10636,WX10639,
    WX10640,WX10645,WX10656,WX10646,WX10652,WX10649,WX10650,WX10653,WX10654,
    WX10659,WX10670,WX10660,WX10666,WX10663,WX10664,WX10667,WX10668,WX10673,
    WX10684,WX10674,WX10680,WX10677,WX10678,WX10681,WX10682,WX10687,WX10698,
    WX10688,WX10694,WX10691,WX10692,WX10695,WX10696,WX10701,WX10712,WX10702,
    WX10708,WX10705,WX10706,WX10709,WX10710,WX10715,WX10726,WX10716,WX10722,
    WX10719,WX10720,WX10723,WX10724,WX10729,WX10740,WX10730,WX10736,WX10733,
    WX10734,WX10737,WX10738,WX10743,WX10754,WX10744,WX10750,WX10747,WX10748,
    WX10751,WX10752,WX10757,WX10768,WX10758,WX10764,WX10761,WX10762,WX10765,
    WX10766,WX10771,WX10782,WX10772,WX10778,WX10775,WX10776,WX10779,WX10780,
    WX10785,WX10796,WX10786,WX10792,WX10789,WX10790,WX10793,WX10794,WX10799,
    WX10810,WX10800,WX10806,WX10803,WX10804,WX10807,WX10808,WX10813,WX10824,
    WX10814,WX10820,WX10817,WX10818,WX10821,WX10822,WX11351,WX11350,WX11352,
    WX11358,WX11357,WX11359,WX11365,WX11364,WX11366,WX11372,WX11371,WX11373,
    WX11379,WX11378,WX11380,WX11386,WX11385,WX11387,WX11393,WX11392,WX11394,
    WX11400,WX11399,WX11401,WX11407,WX11406,WX11408,WX11414,WX11413,WX11415,
    WX11421,WX11420,WX11422,WX11428,WX11427,WX11429,WX11435,WX11434,WX11436,
    WX11442,WX11441,WX11443,WX11449,WX11448,WX11450,WX11456,WX11455,WX11457,
    WX11463,WX11462,WX11464,WX11470,WX11469,WX11471,WX11477,WX11476,WX11478,
    WX11484,WX11483,WX11485,WX11491,WX11490,WX11492,WX11498,WX11497,WX11499,
    WX11505,WX11504,WX11506,WX11512,WX11511,WX11513,WX11519,WX11518,WX11520,
    WX11526,WX11525,WX11527,WX11533,WX11532,WX11534,WX11540,WX11539,WX11541,
    WX11547,WX11546,WX11548,WX11554,WX11553,WX11555,WX11561,WX11560,WX11562,
    WX11568,WX11567,WX11569,WX11578,WX11606,WX11605,WX11604,WX11577,WX11603,
    WX11602,WX11601,WX11600,WX11599,WX11598,WX11576,WX11597,WX11596,WX11595,
    WX11594,WX11575,WX11593,WX11592,WX11591,WX11590,WX11589,WX11588,WX11587,
    WX11586,WX11585,WX11584,WX11583,WX11582,WX11581,WX11580,WX11579,II1988,
    II1989,II1990,II1987,II1995,II1996,II1997,II1986,II2003,II2004,II2005,
    II2002,II2010,II2011,II2012,II2019,II2020,II2021,II2018,II2026,II2027,
    II2028,II2017,II2034,II2035,II2036,II2033,II2041,II2042,II2043,II2050,
    II2051,II2052,II2049,II2057,II2058,II2059,II2048,II2065,II2066,II2067,
    II2064,II2072,II2073,II2074,II2081,II2082,II2083,II2080,II2088,II2089,
    II2090,II2079,II2096,II2097,II2098,II2095,II2103,II2104,II2105,II2112,
    II2113,II2114,II2111,II2119,II2120,II2121,II2110,II2127,II2128,II2129,
    II2126,II2134,II2135,II2136,II2143,II2144,II2145,II2142,II2150,II2151,
    II2152,II2141,II2158,II2159,II2160,II2157,II2165,II2166,II2167,II2174,
    II2175,II2176,II2173,II2181,II2182,II2183,II2172,II2189,II2190,II2191,
    II2188,II2196,II2197,II2198,II2205,II2206,II2207,II2204,II2212,II2213,
    II2214,II2203,II2220,II2221,II2222,II2219,II2227,II2228,II2229,II2236,
    II2237,II2238,II2235,II2243,II2244,II2245,II2234,II2251,II2252,II2253,
    II2250,II2258,II2259,II2260,II2267,II2268,II2269,II2266,II2274,II2275,
    II2276,II2265,II2282,II2283,II2284,II2281,II2289,II2290,II2291,II2298,
    II2299,II2300,II2297,II2305,II2306,II2307,II2296,II2313,II2314,II2315,
    II2312,II2320,II2321,II2322,II2329,II2330,II2331,II2328,II2336,II2337,
    II2338,II2327,II2344,II2345,II2346,II2343,II2351,II2352,II2353,II2360,
    II2361,II2362,II2359,II2367,II2368,II2369,II2358,II2375,II2376,II2377,
    II2374,II2382,II2383,II2384,II2391,II2392,II2393,II2390,II2398,II2399,
    II2400,II2389,II2406,II2407,II2408,II2405,II2413,II2414,II2415,II2422,
    II2423,II2424,II2421,II2429,II2430,II2431,II2420,II2437,II2438,II2439,
    II2436,II2444,II2445,II2446,II2453,II2454,II2455,II2452,II2460,II2461,
    II2462,II2451,II2468,II2469,II2470,II2467,II2475,II2476,II2477,II2484,
    II2485,II2486,II2483,II2491,II2492,II2493,II2482,II2499,II2500,II2501,
    II2498,II2506,II2507,II2508,II2515,II2516,II2517,II2514,II2522,II2523,
    II2524,II2513,II2530,II2531,II2532,II2529,II2537,II2538,II2539,II2546,
    II2547,II2548,II2545,II2553,II2554,II2555,II2544,II2561,II2562,II2563,
    II2560,II2568,II2569,II2570,II2577,II2578,II2579,II2576,II2584,II2585,
    II2586,II2575,II2592,II2593,II2594,II2591,II2599,II2600,II2601,II2608,
    II2609,II2610,II2607,II2615,II2616,II2617,II2606,II2623,II2624,II2625,
    II2622,II2630,II2631,II2632,II2639,II2640,II2641,II2638,II2646,II2647,
    II2648,II2637,II2654,II2655,II2656,II2653,II2661,II2662,II2663,II2670,
    II2671,II2672,II2669,II2677,II2678,II2679,II2668,II2685,II2686,II2687,
    II2684,II2692,II2693,II2694,II2701,II2702,II2703,II2700,II2708,II2709,
    II2710,II2699,II2716,II2717,II2718,II2715,II2723,II2724,II2725,II2732,
    II2733,II2734,II2731,II2739,II2740,II2741,II2730,II2747,II2748,II2749,
    II2746,II2754,II2755,II2756,II2763,II2764,II2765,II2762,II2770,II2771,
    II2772,II2761,II2778,II2779,II2780,II2777,II2785,II2786,II2787,II2794,
    II2795,II2796,II2793,II2801,II2802,II2803,II2792,II2809,II2810,II2811,
    II2808,II2816,II2817,II2818,II2825,II2826,II2827,II2824,II2832,II2833,
    II2834,II2823,II2840,II2841,II2842,II2839,II2847,II2848,II2849,II2856,
    II2857,II2858,II2855,II2863,II2864,II2865,II2854,II2871,II2872,II2873,
    II2870,II2878,II2879,II2880,II2887,II2888,II2889,II2886,II2894,II2895,
    II2896,II2885,II2902,II2903,II2904,II2901,II2909,II2910,II2911,II2918,
    II2919,II2920,II2917,II2925,II2926,II2927,II2916,II2933,II2934,II2935,
    II2932,II2940,II2941,II2942,II2949,II2950,II2951,II2948,II2956,II2957,
    II2958,II2947,II2964,II2965,II2966,II2963,II2971,II2972,II2973,II3052,
    II3053,II3054,II3065,II3066,II3067,II3078,II3079,II3080,II3091,II3092,
    II3093,II3104,II3105,II3106,II3117,II3118,II3119,II3130,II3131,II3132,
    II3143,II3144,II3145,II3156,II3157,II3158,II3169,II3170,II3171,II3182,
    II3183,II3184,II3195,II3196,II3197,II3208,II3209,II3210,II3221,II3222,
    II3223,II3234,II3235,II3236,II3247,II3248,II3249,II3260,II3261,II3262,
    II3273,II3274,II3275,II3286,II3287,II3288,II3299,II3300,II3301,II3312,
    II3313,II3314,II3325,II3326,II3327,II3338,II3339,II3340,II3351,II3352,
    II3353,II3364,II3365,II3366,II3377,II3378,II3379,II3390,II3391,II3392,
    II3403,II3404,II3405,II3416,II3417,II3418,II3429,II3430,II3431,II3442,
    II3443,II3444,II3455,II3456,II3457,II3470,II3471,II3472,II3469,II3477,
    II3478,II3479,II3485,II3486,II3487,II3484,II3492,II3493,II3494,II3500,
    II3501,II3502,II3499,II3507,II3508,II3509,II3514,II3515,II3516,II3521,
    II3522,II3523,II3528,II3529,II3530,II3535,II3536,II3537,II3542,II3543,
    II3544,II3549,II3550,II3551,II3556,II3557,II3558,II3563,II3564,II3565,
    II3570,II3571,II3572,II3577,II3578,II3579,II3584,II3585,II3586,II3591,
    II3592,II3593,II3598,II3599,II3600,II3605,II3606,II3607,II3612,II3613,
    II3614,II3619,II3620,II3621,II3626,II3627,II3628,II3633,II3634,II3635,
    II3640,II3641,II3642,II3647,II3648,II3649,II3654,II3655,II3656,II3661,
    II3662,II3663,II3668,II3669,II3670,II3675,II3676,II3677,II3682,II3683,
    II3684,II3689,II3690,II3691,II3696,II3697,II3698,II3703,II3704,II3705,
    II3710,II3711,II3712,II5993,II5994,II5995,II5992,II6000,II6001,II6002,
    II5991,II6008,II6009,II6010,II6007,II6015,II6016,II6017,II6024,II6025,
    II6026,II6023,II6031,II6032,II6033,II6022,II6039,II6040,II6041,II6038,
    II6046,II6047,II6048,II6055,II6056,II6057,II6054,II6062,II6063,II6064,
    II6053,II6070,II6071,II6072,II6069,II6077,II6078,II6079,II6086,II6087,
    II6088,II6085,II6093,II6094,II6095,II6084,II6101,II6102,II6103,II6100,
    II6108,II6109,II6110,II6117,II6118,II6119,II6116,II6124,II6125,II6126,
    II6115,II6132,II6133,II6134,II6131,II6139,II6140,II6141,II6148,II6149,
    II6150,II6147,II6155,II6156,II6157,II6146,II6163,II6164,II6165,II6162,
    II6170,II6171,II6172,II6179,II6180,II6181,II6178,II6186,II6187,II6188,
    II6177,II6194,II6195,II6196,II6193,II6201,II6202,II6203,II6210,II6211,
    II6212,II6209,II6217,II6218,II6219,II6208,II6225,II6226,II6227,II6224,
    II6232,II6233,II6234,II6241,II6242,II6243,II6240,II6248,II6249,II6250,
    II6239,II6256,II6257,II6258,II6255,II6263,II6264,II6265,II6272,II6273,
    II6274,II6271,II6279,II6280,II6281,II6270,II6287,II6288,II6289,II6286,
    II6294,II6295,II6296,II6303,II6304,II6305,II6302,II6310,II6311,II6312,
    II6301,II6318,II6319,II6320,II6317,II6325,II6326,II6327,II6334,II6335,
    II6336,II6333,II6341,II6342,II6343,II6332,II6349,II6350,II6351,II6348,
    II6356,II6357,II6358,II6365,II6366,II6367,II6364,II6372,II6373,II6374,
    II6363,II6380,II6381,II6382,II6379,II6387,II6388,II6389,II6396,II6397,
    II6398,II6395,II6403,II6404,II6405,II6394,II6411,II6412,II6413,II6410,
    II6418,II6419,II6420,II6427,II6428,II6429,II6426,II6434,II6435,II6436,
    II6425,II6442,II6443,II6444,II6441,II6449,II6450,II6451,II6458,II6459,
    II6460,II6457,II6465,II6466,II6467,II6456,II6473,II6474,II6475,II6472,
    II6480,II6481,II6482,II6489,II6490,II6491,II6488,II6496,II6497,II6498,
    II6487,II6504,II6505,II6506,II6503,II6511,II6512,II6513,II6520,II6521,
    II6522,II6519,II6527,II6528,II6529,II6518,II6535,II6536,II6537,II6534,
    II6542,II6543,II6544,II6551,II6552,II6553,II6550,II6558,II6559,II6560,
    II6549,II6566,II6567,II6568,II6565,II6573,II6574,II6575,II6582,II6583,
    II6584,II6581,II6589,II6590,II6591,II6580,II6597,II6598,II6599,II6596,
    II6604,II6605,II6606,II6613,II6614,II6615,II6612,II6620,II6621,II6622,
    II6611,II6628,II6629,II6630,II6627,II6635,II6636,II6637,II6644,II6645,
    II6646,II6643,II6651,II6652,II6653,II6642,II6659,II6660,II6661,II6658,
    II6666,II6667,II6668,II6675,II6676,II6677,II6674,II6682,II6683,II6684,
    II6673,II6690,II6691,II6692,II6689,II6697,II6698,II6699,II6706,II6707,
    II6708,II6705,II6713,II6714,II6715,II6704,II6721,II6722,II6723,II6720,
    II6728,II6729,II6730,II6737,II6738,II6739,II6736,II6744,II6745,II6746,
    II6735,II6752,II6753,II6754,II6751,II6759,II6760,II6761,II6768,II6769,
    II6770,II6767,II6775,II6776,II6777,II6766,II6783,II6784,II6785,II6782,
    II6790,II6791,II6792,II6799,II6800,II6801,II6798,II6806,II6807,II6808,
    II6797,II6814,II6815,II6816,II6813,II6821,II6822,II6823,II6830,II6831,
    II6832,II6829,II6837,II6838,II6839,II6828,II6845,II6846,II6847,II6844,
    II6852,II6853,II6854,II6861,II6862,II6863,II6860,II6868,II6869,II6870,
    II6859,II6876,II6877,II6878,II6875,II6883,II6884,II6885,II6892,II6893,
    II6894,II6891,II6899,II6900,II6901,II6890,II6907,II6908,II6909,II6906,
    II6914,II6915,II6916,II6923,II6924,II6925,II6922,II6930,II6931,II6932,
    II6921,II6938,II6939,II6940,II6937,II6945,II6946,II6947,II6954,II6955,
    II6956,II6953,II6961,II6962,II6963,II6952,II6969,II6970,II6971,II6968,
    II6976,II6977,II6978,II7057,II7058,II7059,II7070,II7071,II7072,II7083,
    II7084,II7085,II7096,II7097,II7098,II7109,II7110,II7111,II7122,II7123,
    II7124,II7135,II7136,II7137,II7148,II7149,II7150,II7161,II7162,II7163,
    II7174,II7175,II7176,II7187,II7188,II7189,II7200,II7201,II7202,II7213,
    II7214,II7215,II7226,II7227,II7228,II7239,II7240,II7241,II7252,II7253,
    II7254,II7265,II7266,II7267,II7278,II7279,II7280,II7291,II7292,II7293,
    II7304,II7305,II7306,II7317,II7318,II7319,II7330,II7331,II7332,II7343,
    II7344,II7345,II7356,II7357,II7358,II7369,II7370,II7371,II7382,II7383,
    II7384,II7395,II7396,II7397,II7408,II7409,II7410,II7421,II7422,II7423,
    II7434,II7435,II7436,II7447,II7448,II7449,II7460,II7461,II7462,II7475,
    II7476,II7477,II7474,II7482,II7483,II7484,II7490,II7491,II7492,II7489,
    II7497,II7498,II7499,II7505,II7506,II7507,II7504,II7512,II7513,II7514,
    II7519,II7520,II7521,II7526,II7527,II7528,II7533,II7534,II7535,II7540,
    II7541,II7542,II7547,II7548,II7549,II7554,II7555,II7556,II7561,II7562,
    II7563,II7568,II7569,II7570,II7575,II7576,II7577,II7582,II7583,II7584,
    II7589,II7590,II7591,II7596,II7597,II7598,II7603,II7604,II7605,II7610,
    II7611,II7612,II7617,II7618,II7619,II7624,II7625,II7626,II7631,II7632,
    II7633,II7638,II7639,II7640,II7645,II7646,II7647,II7652,II7653,II7654,
    II7659,II7660,II7661,II7666,II7667,II7668,II7673,II7674,II7675,II7680,
    II7681,II7682,II7687,II7688,II7689,II7694,II7695,II7696,II7701,II7702,
    II7703,II7708,II7709,II7710,II7715,II7716,II7717,II9998,II9999,II10000,
    II9997,II10005,II10006,II10007,II9996,II10013,II10014,II10015,II10012,
    II10020,II10021,II10022,II10029,II10030,II10031,II10028,II10036,II10037,
    II10038,II10027,II10044,II10045,II10046,II10043,II10051,II10052,II10053,
    II10060,II10061,II10062,II10059,II10067,II10068,II10069,II10058,II10075,
    II10076,II10077,II10074,II10082,II10083,II10084,II10091,II10092,II10093,
    II10090,II10098,II10099,II10100,II10089,II10106,II10107,II10108,II10105,
    II10113,II10114,II10115,II10122,II10123,II10124,II10121,II10129,II10130,
    II10131,II10120,II10137,II10138,II10139,II10136,II10144,II10145,II10146,
    II10153,II10154,II10155,II10152,II10160,II10161,II10162,II10151,II10168,
    II10169,II10170,II10167,II10175,II10176,II10177,II10184,II10185,II10186,
    II10183,II10191,II10192,II10193,II10182,II10199,II10200,II10201,II10198,
    II10206,II10207,II10208,II10215,II10216,II10217,II10214,II10222,II10223,
    II10224,II10213,II10230,II10231,II10232,II10229,II10237,II10238,II10239,
    II10246,II10247,II10248,II10245,II10253,II10254,II10255,II10244,II10261,
    II10262,II10263,II10260,II10268,II10269,II10270,II10277,II10278,II10279,
    II10276,II10284,II10285,II10286,II10275,II10292,II10293,II10294,II10291,
    II10299,II10300,II10301,II10308,II10309,II10310,II10307,II10315,II10316,
    II10317,II10306,II10323,II10324,II10325,II10322,II10330,II10331,II10332,
    II10339,II10340,II10341,II10338,II10346,II10347,II10348,II10337,II10354,
    II10355,II10356,II10353,II10361,II10362,II10363,II10370,II10371,II10372,
    II10369,II10377,II10378,II10379,II10368,II10385,II10386,II10387,II10384,
    II10392,II10393,II10394,II10401,II10402,II10403,II10400,II10408,II10409,
    II10410,II10399,II10416,II10417,II10418,II10415,II10423,II10424,II10425,
    II10432,II10433,II10434,II10431,II10439,II10440,II10441,II10430,II10447,
    II10448,II10449,II10446,II10454,II10455,II10456,II10463,II10464,II10465,
    II10462,II10470,II10471,II10472,II10461,II10478,II10479,II10480,II10477,
    II10485,II10486,II10487,II10494,II10495,II10496,II10493,II10501,II10502,
    II10503,II10492,II10509,II10510,II10511,II10508,II10516,II10517,II10518,
    II10525,II10526,II10527,II10524,II10532,II10533,II10534,II10523,II10540,
    II10541,II10542,II10539,II10547,II10548,II10549,II10556,II10557,II10558,
    II10555,II10563,II10564,II10565,II10554,II10571,II10572,II10573,II10570,
    II10578,II10579,II10580,II10587,II10588,II10589,II10586,II10594,II10595,
    II10596,II10585,II10602,II10603,II10604,II10601,II10609,II10610,II10611,
    II10618,II10619,II10620,II10617,II10625,II10626,II10627,II10616,II10633,
    II10634,II10635,II10632,II10640,II10641,II10642,II10649,II10650,II10651,
    II10648,II10656,II10657,II10658,II10647,II10664,II10665,II10666,II10663,
    II10671,II10672,II10673,II10680,II10681,II10682,II10679,II10687,II10688,
    II10689,II10678,II10695,II10696,II10697,II10694,II10702,II10703,II10704,
    II10711,II10712,II10713,II10710,II10718,II10719,II10720,II10709,II10726,
    II10727,II10728,II10725,II10733,II10734,II10735,II10742,II10743,II10744,
    II10741,II10749,II10750,II10751,II10740,II10757,II10758,II10759,II10756,
    II10764,II10765,II10766,II10773,II10774,II10775,II10772,II10780,II10781,
    II10782,II10771,II10788,II10789,II10790,II10787,II10795,II10796,II10797,
    II10804,II10805,II10806,II10803,II10811,II10812,II10813,II10802,II10819,
    II10820,II10821,II10818,II10826,II10827,II10828,II10835,II10836,II10837,
    II10834,II10842,II10843,II10844,II10833,II10850,II10851,II10852,II10849,
    II10857,II10858,II10859,II10866,II10867,II10868,II10865,II10873,II10874,
    II10875,II10864,II10881,II10882,II10883,II10880,II10888,II10889,II10890,
    II10897,II10898,II10899,II10896,II10904,II10905,II10906,II10895,II10912,
    II10913,II10914,II10911,II10919,II10920,II10921,II10928,II10929,II10930,
    II10927,II10935,II10936,II10937,II10926,II10943,II10944,II10945,II10942,
    II10950,II10951,II10952,II10959,II10960,II10961,II10958,II10966,II10967,
    II10968,II10957,II10974,II10975,II10976,II10973,II10981,II10982,II10983,
    II11062,II11063,II11064,II11075,II11076,II11077,II11088,II11089,II11090,
    II11101,II11102,II11103,II11114,II11115,II11116,II11127,II11128,II11129,
    II11140,II11141,II11142,II11153,II11154,II11155,II11166,II11167,II11168,
    II11179,II11180,II11181,II11192,II11193,II11194,II11205,II11206,II11207,
    II11218,II11219,II11220,II11231,II11232,II11233,II11244,II11245,II11246,
    II11257,II11258,II11259,II11270,II11271,II11272,II11283,II11284,II11285,
    II11296,II11297,II11298,II11309,II11310,II11311,II11322,II11323,II11324,
    II11335,II11336,II11337,II11348,II11349,II11350,II11361,II11362,II11363,
    II11374,II11375,II11376,II11387,II11388,II11389,II11400,II11401,II11402,
    II11413,II11414,II11415,II11426,II11427,II11428,II11439,II11440,II11441,
    II11452,II11453,II11454,II11465,II11466,II11467,II11480,II11481,II11482,
    II11479,II11487,II11488,II11489,II11495,II11496,II11497,II11494,II11502,
    II11503,II11504,II11510,II11511,II11512,II11509,II11517,II11518,II11519,
    II11524,II11525,II11526,II11531,II11532,II11533,II11538,II11539,II11540,
    II11545,II11546,II11547,II11552,II11553,II11554,II11559,II11560,II11561,
    II11566,II11567,II11568,II11573,II11574,II11575,II11580,II11581,II11582,
    II11587,II11588,II11589,II11594,II11595,II11596,II11601,II11602,II11603,
    II11608,II11609,II11610,II11615,II11616,II11617,II11622,II11623,II11624,
    II11629,II11630,II11631,II11636,II11637,II11638,II11643,II11644,II11645,
    II11650,II11651,II11652,II11657,II11658,II11659,II11664,II11665,II11666,
    II11671,II11672,II11673,II11678,II11679,II11680,II11685,II11686,II11687,
    II11692,II11693,II11694,II11699,II11700,II11701,II11706,II11707,II11708,
    II11713,II11714,II11715,II11720,II11721,II11722,II14003,II14004,II14005,
    II14002,II14010,II14011,II14012,II14001,II14018,II14019,II14020,II14017,
    II14025,II14026,II14027,II14034,II14035,II14036,II14033,II14041,II14042,
    II14043,II14032,II14049,II14050,II14051,II14048,II14056,II14057,II14058,
    II14065,II14066,II14067,II14064,II14072,II14073,II14074,II14063,II14080,
    II14081,II14082,II14079,II14087,II14088,II14089,II14096,II14097,II14098,
    II14095,II14103,II14104,II14105,II14094,II14111,II14112,II14113,II14110,
    II14118,II14119,II14120,II14127,II14128,II14129,II14126,II14134,II14135,
    II14136,II14125,II14142,II14143,II14144,II14141,II14149,II14150,II14151,
    II14158,II14159,II14160,II14157,II14165,II14166,II14167,II14156,II14173,
    II14174,II14175,II14172,II14180,II14181,II14182,II14189,II14190,II14191,
    II14188,II14196,II14197,II14198,II14187,II14204,II14205,II14206,II14203,
    II14211,II14212,II14213,II14220,II14221,II14222,II14219,II14227,II14228,
    II14229,II14218,II14235,II14236,II14237,II14234,II14242,II14243,II14244,
    II14251,II14252,II14253,II14250,II14258,II14259,II14260,II14249,II14266,
    II14267,II14268,II14265,II14273,II14274,II14275,II14282,II14283,II14284,
    II14281,II14289,II14290,II14291,II14280,II14297,II14298,II14299,II14296,
    II14304,II14305,II14306,II14313,II14314,II14315,II14312,II14320,II14321,
    II14322,II14311,II14328,II14329,II14330,II14327,II14335,II14336,II14337,
    II14344,II14345,II14346,II14343,II14351,II14352,II14353,II14342,II14359,
    II14360,II14361,II14358,II14366,II14367,II14368,II14375,II14376,II14377,
    II14374,II14382,II14383,II14384,II14373,II14390,II14391,II14392,II14389,
    II14397,II14398,II14399,II14406,II14407,II14408,II14405,II14413,II14414,
    II14415,II14404,II14421,II14422,II14423,II14420,II14428,II14429,II14430,
    II14437,II14438,II14439,II14436,II14444,II14445,II14446,II14435,II14452,
    II14453,II14454,II14451,II14459,II14460,II14461,II14468,II14469,II14470,
    II14467,II14475,II14476,II14477,II14466,II14483,II14484,II14485,II14482,
    II14490,II14491,II14492,II14499,II14500,II14501,II14498,II14506,II14507,
    II14508,II14497,II14514,II14515,II14516,II14513,II14521,II14522,II14523,
    II14530,II14531,II14532,II14529,II14537,II14538,II14539,II14528,II14545,
    II14546,II14547,II14544,II14552,II14553,II14554,II14561,II14562,II14563,
    II14560,II14568,II14569,II14570,II14559,II14576,II14577,II14578,II14575,
    II14583,II14584,II14585,II14592,II14593,II14594,II14591,II14599,II14600,
    II14601,II14590,II14607,II14608,II14609,II14606,II14614,II14615,II14616,
    II14623,II14624,II14625,II14622,II14630,II14631,II14632,II14621,II14638,
    II14639,II14640,II14637,II14645,II14646,II14647,II14654,II14655,II14656,
    II14653,II14661,II14662,II14663,II14652,II14669,II14670,II14671,II14668,
    II14676,II14677,II14678,II14685,II14686,II14687,II14684,II14692,II14693,
    II14694,II14683,II14700,II14701,II14702,II14699,II14707,II14708,II14709,
    II14716,II14717,II14718,II14715,II14723,II14724,II14725,II14714,II14731,
    II14732,II14733,II14730,II14738,II14739,II14740,II14747,II14748,II14749,
    II14746,II14754,II14755,II14756,II14745,II14762,II14763,II14764,II14761,
    II14769,II14770,II14771,II14778,II14779,II14780,II14777,II14785,II14786,
    II14787,II14776,II14793,II14794,II14795,II14792,II14800,II14801,II14802,
    II14809,II14810,II14811,II14808,II14816,II14817,II14818,II14807,II14824,
    II14825,II14826,II14823,II14831,II14832,II14833,II14840,II14841,II14842,
    II14839,II14847,II14848,II14849,II14838,II14855,II14856,II14857,II14854,
    II14862,II14863,II14864,II14871,II14872,II14873,II14870,II14878,II14879,
    II14880,II14869,II14886,II14887,II14888,II14885,II14893,II14894,II14895,
    II14902,II14903,II14904,II14901,II14909,II14910,II14911,II14900,II14917,
    II14918,II14919,II14916,II14924,II14925,II14926,II14933,II14934,II14935,
    II14932,II14940,II14941,II14942,II14931,II14948,II14949,II14950,II14947,
    II14955,II14956,II14957,II14964,II14965,II14966,II14963,II14971,II14972,
    II14973,II14962,II14979,II14980,II14981,II14978,II14986,II14987,II14988,
    II15067,II15068,II15069,II15080,II15081,II15082,II15093,II15094,II15095,
    II15106,II15107,II15108,II15119,II15120,II15121,II15132,II15133,II15134,
    II15145,II15146,II15147,II15158,II15159,II15160,II15171,II15172,II15173,
    II15184,II15185,II15186,II15197,II15198,II15199,II15210,II15211,II15212,
    II15223,II15224,II15225,II15236,II15237,II15238,II15249,II15250,II15251,
    II15262,II15263,II15264,II15275,II15276,II15277,II15288,II15289,II15290,
    II15301,II15302,II15303,II15314,II15315,II15316,II15327,II15328,II15329,
    II15340,II15341,II15342,II15353,II15354,II15355,II15366,II15367,II15368,
    II15379,II15380,II15381,II15392,II15393,II15394,II15405,II15406,II15407,
    II15418,II15419,II15420,II15431,II15432,II15433,II15444,II15445,II15446,
    II15457,II15458,II15459,II15470,II15471,II15472,II15485,II15486,II15487,
    II15484,II15492,II15493,II15494,II15500,II15501,II15502,II15499,II15507,
    II15508,II15509,II15515,II15516,II15517,II15514,II15522,II15523,II15524,
    II15529,II15530,II15531,II15536,II15537,II15538,II15543,II15544,II15545,
    II15550,II15551,II15552,II15557,II15558,II15559,II15564,II15565,II15566,
    II15571,II15572,II15573,II15578,II15579,II15580,II15585,II15586,II15587,
    II15592,II15593,II15594,II15599,II15600,II15601,II15606,II15607,II15608,
    II15613,II15614,II15615,II15620,II15621,II15622,II15627,II15628,II15629,
    II15634,II15635,II15636,II15641,II15642,II15643,II15648,II15649,II15650,
    II15655,II15656,II15657,II15662,II15663,II15664,II15669,II15670,II15671,
    II15676,II15677,II15678,II15683,II15684,II15685,II15690,II15691,II15692,
    II15697,II15698,II15699,II15704,II15705,II15706,II15711,II15712,II15713,
    II15718,II15719,II15720,II15725,II15726,II15727,II18008,II18009,II18010,
    II18007,II18015,II18016,II18017,II18006,II18023,II18024,II18025,II18022,
    II18030,II18031,II18032,II18039,II18040,II18041,II18038,II18046,II18047,
    II18048,II18037,II18054,II18055,II18056,II18053,II18061,II18062,II18063,
    II18070,II18071,II18072,II18069,II18077,II18078,II18079,II18068,II18085,
    II18086,II18087,II18084,II18092,II18093,II18094,II18101,II18102,II18103,
    II18100,II18108,II18109,II18110,II18099,II18116,II18117,II18118,II18115,
    II18123,II18124,II18125,II18132,II18133,II18134,II18131,II18139,II18140,
    II18141,II18130,II18147,II18148,II18149,II18146,II18154,II18155,II18156,
    II18163,II18164,II18165,II18162,II18170,II18171,II18172,II18161,II18178,
    II18179,II18180,II18177,II18185,II18186,II18187,II18194,II18195,II18196,
    II18193,II18201,II18202,II18203,II18192,II18209,II18210,II18211,II18208,
    II18216,II18217,II18218,II18225,II18226,II18227,II18224,II18232,II18233,
    II18234,II18223,II18240,II18241,II18242,II18239,II18247,II18248,II18249,
    II18256,II18257,II18258,II18255,II18263,II18264,II18265,II18254,II18271,
    II18272,II18273,II18270,II18278,II18279,II18280,II18287,II18288,II18289,
    II18286,II18294,II18295,II18296,II18285,II18302,II18303,II18304,II18301,
    II18309,II18310,II18311,II18318,II18319,II18320,II18317,II18325,II18326,
    II18327,II18316,II18333,II18334,II18335,II18332,II18340,II18341,II18342,
    II18349,II18350,II18351,II18348,II18356,II18357,II18358,II18347,II18364,
    II18365,II18366,II18363,II18371,II18372,II18373,II18380,II18381,II18382,
    II18379,II18387,II18388,II18389,II18378,II18395,II18396,II18397,II18394,
    II18402,II18403,II18404,II18411,II18412,II18413,II18410,II18418,II18419,
    II18420,II18409,II18426,II18427,II18428,II18425,II18433,II18434,II18435,
    II18442,II18443,II18444,II18441,II18449,II18450,II18451,II18440,II18457,
    II18458,II18459,II18456,II18464,II18465,II18466,II18473,II18474,II18475,
    II18472,II18480,II18481,II18482,II18471,II18488,II18489,II18490,II18487,
    II18495,II18496,II18497,II18504,II18505,II18506,II18503,II18511,II18512,
    II18513,II18502,II18519,II18520,II18521,II18518,II18526,II18527,II18528,
    II18535,II18536,II18537,II18534,II18542,II18543,II18544,II18533,II18550,
    II18551,II18552,II18549,II18557,II18558,II18559,II18566,II18567,II18568,
    II18565,II18573,II18574,II18575,II18564,II18581,II18582,II18583,II18580,
    II18588,II18589,II18590,II18597,II18598,II18599,II18596,II18604,II18605,
    II18606,II18595,II18612,II18613,II18614,II18611,II18619,II18620,II18621,
    II18628,II18629,II18630,II18627,II18635,II18636,II18637,II18626,II18643,
    II18644,II18645,II18642,II18650,II18651,II18652,II18659,II18660,II18661,
    II18658,II18666,II18667,II18668,II18657,II18674,II18675,II18676,II18673,
    II18681,II18682,II18683,II18690,II18691,II18692,II18689,II18697,II18698,
    II18699,II18688,II18705,II18706,II18707,II18704,II18712,II18713,II18714,
    II18721,II18722,II18723,II18720,II18728,II18729,II18730,II18719,II18736,
    II18737,II18738,II18735,II18743,II18744,II18745,II18752,II18753,II18754,
    II18751,II18759,II18760,II18761,II18750,II18767,II18768,II18769,II18766,
    II18774,II18775,II18776,II18783,II18784,II18785,II18782,II18790,II18791,
    II18792,II18781,II18798,II18799,II18800,II18797,II18805,II18806,II18807,
    II18814,II18815,II18816,II18813,II18821,II18822,II18823,II18812,II18829,
    II18830,II18831,II18828,II18836,II18837,II18838,II18845,II18846,II18847,
    II18844,II18852,II18853,II18854,II18843,II18860,II18861,II18862,II18859,
    II18867,II18868,II18869,II18876,II18877,II18878,II18875,II18883,II18884,
    II18885,II18874,II18891,II18892,II18893,II18890,II18898,II18899,II18900,
    II18907,II18908,II18909,II18906,II18914,II18915,II18916,II18905,II18922,
    II18923,II18924,II18921,II18929,II18930,II18931,II18938,II18939,II18940,
    II18937,II18945,II18946,II18947,II18936,II18953,II18954,II18955,II18952,
    II18960,II18961,II18962,II18969,II18970,II18971,II18968,II18976,II18977,
    II18978,II18967,II18984,II18985,II18986,II18983,II18991,II18992,II18993,
    II19072,II19073,II19074,II19085,II19086,II19087,II19098,II19099,II19100,
    II19111,II19112,II19113,II19124,II19125,II19126,II19137,II19138,II19139,
    II19150,II19151,II19152,II19163,II19164,II19165,II19176,II19177,II19178,
    II19189,II19190,II19191,II19202,II19203,II19204,II19215,II19216,II19217,
    II19228,II19229,II19230,II19241,II19242,II19243,II19254,II19255,II19256,
    II19267,II19268,II19269,II19280,II19281,II19282,II19293,II19294,II19295,
    II19306,II19307,II19308,II19319,II19320,II19321,II19332,II19333,II19334,
    II19345,II19346,II19347,II19358,II19359,II19360,II19371,II19372,II19373,
    II19384,II19385,II19386,II19397,II19398,II19399,II19410,II19411,II19412,
    II19423,II19424,II19425,II19436,II19437,II19438,II19449,II19450,II19451,
    II19462,II19463,II19464,II19475,II19476,II19477,II19490,II19491,II19492,
    II19489,II19497,II19498,II19499,II19505,II19506,II19507,II19504,II19512,
    II19513,II19514,II19520,II19521,II19522,II19519,II19527,II19528,II19529,
    II19534,II19535,II19536,II19541,II19542,II19543,II19548,II19549,II19550,
    II19555,II19556,II19557,II19562,II19563,II19564,II19569,II19570,II19571,
    II19576,II19577,II19578,II19583,II19584,II19585,II19590,II19591,II19592,
    II19597,II19598,II19599,II19604,II19605,II19606,II19611,II19612,II19613,
    II19618,II19619,II19620,II19625,II19626,II19627,II19632,II19633,II19634,
    II19639,II19640,II19641,II19646,II19647,II19648,II19653,II19654,II19655,
    II19660,II19661,II19662,II19667,II19668,II19669,II19674,II19675,II19676,
    II19681,II19682,II19683,II19688,II19689,II19690,II19695,II19696,II19697,
    II19702,II19703,II19704,II19709,II19710,II19711,II19716,II19717,II19718,
    II19723,II19724,II19725,II19730,II19731,II19732,II22013,II22014,II22015,
    II22012,II22020,II22021,II22022,II22011,II22028,II22029,II22030,II22027,
    II22035,II22036,II22037,II22044,II22045,II22046,II22043,II22051,II22052,
    II22053,II22042,II22059,II22060,II22061,II22058,II22066,II22067,II22068,
    II22075,II22076,II22077,II22074,II22082,II22083,II22084,II22073,II22090,
    II22091,II22092,II22089,II22097,II22098,II22099,II22106,II22107,II22108,
    II22105,II22113,II22114,II22115,II22104,II22121,II22122,II22123,II22120,
    II22128,II22129,II22130,II22137,II22138,II22139,II22136,II22144,II22145,
    II22146,II22135,II22152,II22153,II22154,II22151,II22159,II22160,II22161,
    II22168,II22169,II22170,II22167,II22175,II22176,II22177,II22166,II22183,
    II22184,II22185,II22182,II22190,II22191,II22192,II22199,II22200,II22201,
    II22198,II22206,II22207,II22208,II22197,II22214,II22215,II22216,II22213,
    II22221,II22222,II22223,II22230,II22231,II22232,II22229,II22237,II22238,
    II22239,II22228,II22245,II22246,II22247,II22244,II22252,II22253,II22254,
    II22261,II22262,II22263,II22260,II22268,II22269,II22270,II22259,II22276,
    II22277,II22278,II22275,II22283,II22284,II22285,II22292,II22293,II22294,
    II22291,II22299,II22300,II22301,II22290,II22307,II22308,II22309,II22306,
    II22314,II22315,II22316,II22323,II22324,II22325,II22322,II22330,II22331,
    II22332,II22321,II22338,II22339,II22340,II22337,II22345,II22346,II22347,
    II22354,II22355,II22356,II22353,II22361,II22362,II22363,II22352,II22369,
    II22370,II22371,II22368,II22376,II22377,II22378,II22385,II22386,II22387,
    II22384,II22392,II22393,II22394,II22383,II22400,II22401,II22402,II22399,
    II22407,II22408,II22409,II22416,II22417,II22418,II22415,II22423,II22424,
    II22425,II22414,II22431,II22432,II22433,II22430,II22438,II22439,II22440,
    II22447,II22448,II22449,II22446,II22454,II22455,II22456,II22445,II22462,
    II22463,II22464,II22461,II22469,II22470,II22471,II22478,II22479,II22480,
    II22477,II22485,II22486,II22487,II22476,II22493,II22494,II22495,II22492,
    II22500,II22501,II22502,II22509,II22510,II22511,II22508,II22516,II22517,
    II22518,II22507,II22524,II22525,II22526,II22523,II22531,II22532,II22533,
    II22540,II22541,II22542,II22539,II22547,II22548,II22549,II22538,II22555,
    II22556,II22557,II22554,II22562,II22563,II22564,II22571,II22572,II22573,
    II22570,II22578,II22579,II22580,II22569,II22586,II22587,II22588,II22585,
    II22593,II22594,II22595,II22602,II22603,II22604,II22601,II22609,II22610,
    II22611,II22600,II22617,II22618,II22619,II22616,II22624,II22625,II22626,
    II22633,II22634,II22635,II22632,II22640,II22641,II22642,II22631,II22648,
    II22649,II22650,II22647,II22655,II22656,II22657,II22664,II22665,II22666,
    II22663,II22671,II22672,II22673,II22662,II22679,II22680,II22681,II22678,
    II22686,II22687,II22688,II22695,II22696,II22697,II22694,II22702,II22703,
    II22704,II22693,II22710,II22711,II22712,II22709,II22717,II22718,II22719,
    II22726,II22727,II22728,II22725,II22733,II22734,II22735,II22724,II22741,
    II22742,II22743,II22740,II22748,II22749,II22750,II22757,II22758,II22759,
    II22756,II22764,II22765,II22766,II22755,II22772,II22773,II22774,II22771,
    II22779,II22780,II22781,II22788,II22789,II22790,II22787,II22795,II22796,
    II22797,II22786,II22803,II22804,II22805,II22802,II22810,II22811,II22812,
    II22819,II22820,II22821,II22818,II22826,II22827,II22828,II22817,II22834,
    II22835,II22836,II22833,II22841,II22842,II22843,II22850,II22851,II22852,
    II22849,II22857,II22858,II22859,II22848,II22865,II22866,II22867,II22864,
    II22872,II22873,II22874,II22881,II22882,II22883,II22880,II22888,II22889,
    II22890,II22879,II22896,II22897,II22898,II22895,II22903,II22904,II22905,
    II22912,II22913,II22914,II22911,II22919,II22920,II22921,II22910,II22927,
    II22928,II22929,II22926,II22934,II22935,II22936,II22943,II22944,II22945,
    II22942,II22950,II22951,II22952,II22941,II22958,II22959,II22960,II22957,
    II22965,II22966,II22967,II22974,II22975,II22976,II22973,II22981,II22982,
    II22983,II22972,II22989,II22990,II22991,II22988,II22996,II22997,II22998,
    II23077,II23078,II23079,II23090,II23091,II23092,II23103,II23104,II23105,
    II23116,II23117,II23118,II23129,II23130,II23131,II23142,II23143,II23144,
    II23155,II23156,II23157,II23168,II23169,II23170,II23181,II23182,II23183,
    II23194,II23195,II23196,II23207,II23208,II23209,II23220,II23221,II23222,
    II23233,II23234,II23235,II23246,II23247,II23248,II23259,II23260,II23261,
    II23272,II23273,II23274,II23285,II23286,II23287,II23298,II23299,II23300,
    II23311,II23312,II23313,II23324,II23325,II23326,II23337,II23338,II23339,
    II23350,II23351,II23352,II23363,II23364,II23365,II23376,II23377,II23378,
    II23389,II23390,II23391,II23402,II23403,II23404,II23415,II23416,II23417,
    II23428,II23429,II23430,II23441,II23442,II23443,II23454,II23455,II23456,
    II23467,II23468,II23469,II23480,II23481,II23482,II23495,II23496,II23497,
    II23494,II23502,II23503,II23504,II23510,II23511,II23512,II23509,II23517,
    II23518,II23519,II23525,II23526,II23527,II23524,II23532,II23533,II23534,
    II23539,II23540,II23541,II23546,II23547,II23548,II23553,II23554,II23555,
    II23560,II23561,II23562,II23567,II23568,II23569,II23574,II23575,II23576,
    II23581,II23582,II23583,II23588,II23589,II23590,II23595,II23596,II23597,
    II23602,II23603,II23604,II23609,II23610,II23611,II23616,II23617,II23618,
    II23623,II23624,II23625,II23630,II23631,II23632,II23637,II23638,II23639,
    II23644,II23645,II23646,II23651,II23652,II23653,II23658,II23659,II23660,
    II23665,II23666,II23667,II23672,II23673,II23674,II23679,II23680,II23681,
    II23686,II23687,II23688,II23693,II23694,II23695,II23700,II23701,II23702,
    II23707,II23708,II23709,II23714,II23715,II23716,II23721,II23722,II23723,
    II23728,II23729,II23730,II23735,II23736,II23737,II26018,II26019,II26020,
    II26017,II26025,II26026,II26027,II26016,II26033,II26034,II26035,II26032,
    II26040,II26041,II26042,II26049,II26050,II26051,II26048,II26056,II26057,
    II26058,II26047,II26064,II26065,II26066,II26063,II26071,II26072,II26073,
    II26080,II26081,II26082,II26079,II26087,II26088,II26089,II26078,II26095,
    II26096,II26097,II26094,II26102,II26103,II26104,II26111,II26112,II26113,
    II26110,II26118,II26119,II26120,II26109,II26126,II26127,II26128,II26125,
    II26133,II26134,II26135,II26142,II26143,II26144,II26141,II26149,II26150,
    II26151,II26140,II26157,II26158,II26159,II26156,II26164,II26165,II26166,
    II26173,II26174,II26175,II26172,II26180,II26181,II26182,II26171,II26188,
    II26189,II26190,II26187,II26195,II26196,II26197,II26204,II26205,II26206,
    II26203,II26211,II26212,II26213,II26202,II26219,II26220,II26221,II26218,
    II26226,II26227,II26228,II26235,II26236,II26237,II26234,II26242,II26243,
    II26244,II26233,II26250,II26251,II26252,II26249,II26257,II26258,II26259,
    II26266,II26267,II26268,II26265,II26273,II26274,II26275,II26264,II26281,
    II26282,II26283,II26280,II26288,II26289,II26290,II26297,II26298,II26299,
    II26296,II26304,II26305,II26306,II26295,II26312,II26313,II26314,II26311,
    II26319,II26320,II26321,II26328,II26329,II26330,II26327,II26335,II26336,
    II26337,II26326,II26343,II26344,II26345,II26342,II26350,II26351,II26352,
    II26359,II26360,II26361,II26358,II26366,II26367,II26368,II26357,II26374,
    II26375,II26376,II26373,II26381,II26382,II26383,II26390,II26391,II26392,
    II26389,II26397,II26398,II26399,II26388,II26405,II26406,II26407,II26404,
    II26412,II26413,II26414,II26421,II26422,II26423,II26420,II26428,II26429,
    II26430,II26419,II26436,II26437,II26438,II26435,II26443,II26444,II26445,
    II26452,II26453,II26454,II26451,II26459,II26460,II26461,II26450,II26467,
    II26468,II26469,II26466,II26474,II26475,II26476,II26483,II26484,II26485,
    II26482,II26490,II26491,II26492,II26481,II26498,II26499,II26500,II26497,
    II26505,II26506,II26507,II26514,II26515,II26516,II26513,II26521,II26522,
    II26523,II26512,II26529,II26530,II26531,II26528,II26536,II26537,II26538,
    II26545,II26546,II26547,II26544,II26552,II26553,II26554,II26543,II26560,
    II26561,II26562,II26559,II26567,II26568,II26569,II26576,II26577,II26578,
    II26575,II26583,II26584,II26585,II26574,II26591,II26592,II26593,II26590,
    II26598,II26599,II26600,II26607,II26608,II26609,II26606,II26614,II26615,
    II26616,II26605,II26622,II26623,II26624,II26621,II26629,II26630,II26631,
    II26638,II26639,II26640,II26637,II26645,II26646,II26647,II26636,II26653,
    II26654,II26655,II26652,II26660,II26661,II26662,II26669,II26670,II26671,
    II26668,II26676,II26677,II26678,II26667,II26684,II26685,II26686,II26683,
    II26691,II26692,II26693,II26700,II26701,II26702,II26699,II26707,II26708,
    II26709,II26698,II26715,II26716,II26717,II26714,II26722,II26723,II26724,
    II26731,II26732,II26733,II26730,II26738,II26739,II26740,II26729,II26746,
    II26747,II26748,II26745,II26753,II26754,II26755,II26762,II26763,II26764,
    II26761,II26769,II26770,II26771,II26760,II26777,II26778,II26779,II26776,
    II26784,II26785,II26786,II26793,II26794,II26795,II26792,II26800,II26801,
    II26802,II26791,II26808,II26809,II26810,II26807,II26815,II26816,II26817,
    II26824,II26825,II26826,II26823,II26831,II26832,II26833,II26822,II26839,
    II26840,II26841,II26838,II26846,II26847,II26848,II26855,II26856,II26857,
    II26854,II26862,II26863,II26864,II26853,II26870,II26871,II26872,II26869,
    II26877,II26878,II26879,II26886,II26887,II26888,II26885,II26893,II26894,
    II26895,II26884,II26901,II26902,II26903,II26900,II26908,II26909,II26910,
    II26917,II26918,II26919,II26916,II26924,II26925,II26926,II26915,II26932,
    II26933,II26934,II26931,II26939,II26940,II26941,II26948,II26949,II26950,
    II26947,II26955,II26956,II26957,II26946,II26963,II26964,II26965,II26962,
    II26970,II26971,II26972,II26979,II26980,II26981,II26978,II26986,II26987,
    II26988,II26977,II26994,II26995,II26996,II26993,II27001,II27002,II27003,
    II27082,II27083,II27084,II27095,II27096,II27097,II27108,II27109,II27110,
    II27121,II27122,II27123,II27134,II27135,II27136,II27147,II27148,II27149,
    II27160,II27161,II27162,II27173,II27174,II27175,II27186,II27187,II27188,
    II27199,II27200,II27201,II27212,II27213,II27214,II27225,II27226,II27227,
    II27238,II27239,II27240,II27251,II27252,II27253,II27264,II27265,II27266,
    II27277,II27278,II27279,II27290,II27291,II27292,II27303,II27304,II27305,
    II27316,II27317,II27318,II27329,II27330,II27331,II27342,II27343,II27344,
    II27355,II27356,II27357,II27368,II27369,II27370,II27381,II27382,II27383,
    II27394,II27395,II27396,II27407,II27408,II27409,II27420,II27421,II27422,
    II27433,II27434,II27435,II27446,II27447,II27448,II27459,II27460,II27461,
    II27472,II27473,II27474,II27485,II27486,II27487,II27500,II27501,II27502,
    II27499,II27507,II27508,II27509,II27515,II27516,II27517,II27514,II27522,
    II27523,II27524,II27530,II27531,II27532,II27529,II27537,II27538,II27539,
    II27544,II27545,II27546,II27551,II27552,II27553,II27558,II27559,II27560,
    II27565,II27566,II27567,II27572,II27573,II27574,II27579,II27580,II27581,
    II27586,II27587,II27588,II27593,II27594,II27595,II27600,II27601,II27602,
    II27607,II27608,II27609,II27614,II27615,II27616,II27621,II27622,II27623,
    II27628,II27629,II27630,II27635,II27636,II27637,II27642,II27643,II27644,
    II27649,II27650,II27651,II27656,II27657,II27658,II27663,II27664,II27665,
    II27670,II27671,II27672,II27677,II27678,II27679,II27684,II27685,II27686,
    II27691,II27692,II27693,II27698,II27699,II27700,II27705,II27706,II27707,
    II27712,II27713,II27714,II27719,II27720,II27721,II27726,II27727,II27728,
    II27733,II27734,II27735,II27740,II27741,II27742,II30023,II30024,II30025,
    II30022,II30030,II30031,II30032,II30021,II30038,II30039,II30040,II30037,
    II30045,II30046,II30047,II30054,II30055,II30056,II30053,II30061,II30062,
    II30063,II30052,II30069,II30070,II30071,II30068,II30076,II30077,II30078,
    II30085,II30086,II30087,II30084,II30092,II30093,II30094,II30083,II30100,
    II30101,II30102,II30099,II30107,II30108,II30109,II30116,II30117,II30118,
    II30115,II30123,II30124,II30125,II30114,II30131,II30132,II30133,II30130,
    II30138,II30139,II30140,II30147,II30148,II30149,II30146,II30154,II30155,
    II30156,II30145,II30162,II30163,II30164,II30161,II30169,II30170,II30171,
    II30178,II30179,II30180,II30177,II30185,II30186,II30187,II30176,II30193,
    II30194,II30195,II30192,II30200,II30201,II30202,II30209,II30210,II30211,
    II30208,II30216,II30217,II30218,II30207,II30224,II30225,II30226,II30223,
    II30231,II30232,II30233,II30240,II30241,II30242,II30239,II30247,II30248,
    II30249,II30238,II30255,II30256,II30257,II30254,II30262,II30263,II30264,
    II30271,II30272,II30273,II30270,II30278,II30279,II30280,II30269,II30286,
    II30287,II30288,II30285,II30293,II30294,II30295,II30302,II30303,II30304,
    II30301,II30309,II30310,II30311,II30300,II30317,II30318,II30319,II30316,
    II30324,II30325,II30326,II30333,II30334,II30335,II30332,II30340,II30341,
    II30342,II30331,II30348,II30349,II30350,II30347,II30355,II30356,II30357,
    II30364,II30365,II30366,II30363,II30371,II30372,II30373,II30362,II30379,
    II30380,II30381,II30378,II30386,II30387,II30388,II30395,II30396,II30397,
    II30394,II30402,II30403,II30404,II30393,II30410,II30411,II30412,II30409,
    II30417,II30418,II30419,II30426,II30427,II30428,II30425,II30433,II30434,
    II30435,II30424,II30441,II30442,II30443,II30440,II30448,II30449,II30450,
    II30457,II30458,II30459,II30456,II30464,II30465,II30466,II30455,II30472,
    II30473,II30474,II30471,II30479,II30480,II30481,II30488,II30489,II30490,
    II30487,II30495,II30496,II30497,II30486,II30503,II30504,II30505,II30502,
    II30510,II30511,II30512,II30519,II30520,II30521,II30518,II30526,II30527,
    II30528,II30517,II30534,II30535,II30536,II30533,II30541,II30542,II30543,
    II30550,II30551,II30552,II30549,II30557,II30558,II30559,II30548,II30565,
    II30566,II30567,II30564,II30572,II30573,II30574,II30581,II30582,II30583,
    II30580,II30588,II30589,II30590,II30579,II30596,II30597,II30598,II30595,
    II30603,II30604,II30605,II30612,II30613,II30614,II30611,II30619,II30620,
    II30621,II30610,II30627,II30628,II30629,II30626,II30634,II30635,II30636,
    II30643,II30644,II30645,II30642,II30650,II30651,II30652,II30641,II30658,
    II30659,II30660,II30657,II30665,II30666,II30667,II30674,II30675,II30676,
    II30673,II30681,II30682,II30683,II30672,II30689,II30690,II30691,II30688,
    II30696,II30697,II30698,II30705,II30706,II30707,II30704,II30712,II30713,
    II30714,II30703,II30720,II30721,II30722,II30719,II30727,II30728,II30729,
    II30736,II30737,II30738,II30735,II30743,II30744,II30745,II30734,II30751,
    II30752,II30753,II30750,II30758,II30759,II30760,II30767,II30768,II30769,
    II30766,II30774,II30775,II30776,II30765,II30782,II30783,II30784,II30781,
    II30789,II30790,II30791,II30798,II30799,II30800,II30797,II30805,II30806,
    II30807,II30796,II30813,II30814,II30815,II30812,II30820,II30821,II30822,
    II30829,II30830,II30831,II30828,II30836,II30837,II30838,II30827,II30844,
    II30845,II30846,II30843,II30851,II30852,II30853,II30860,II30861,II30862,
    II30859,II30867,II30868,II30869,II30858,II30875,II30876,II30877,II30874,
    II30882,II30883,II30884,II30891,II30892,II30893,II30890,II30898,II30899,
    II30900,II30889,II30906,II30907,II30908,II30905,II30913,II30914,II30915,
    II30922,II30923,II30924,II30921,II30929,II30930,II30931,II30920,II30937,
    II30938,II30939,II30936,II30944,II30945,II30946,II30953,II30954,II30955,
    II30952,II30960,II30961,II30962,II30951,II30968,II30969,II30970,II30967,
    II30975,II30976,II30977,II30984,II30985,II30986,II30983,II30991,II30992,
    II30993,II30982,II30999,II31000,II31001,II30998,II31006,II31007,II31008,
    II31087,II31088,II31089,II31100,II31101,II31102,II31113,II31114,II31115,
    II31126,II31127,II31128,II31139,II31140,II31141,II31152,II31153,II31154,
    II31165,II31166,II31167,II31178,II31179,II31180,II31191,II31192,II31193,
    II31204,II31205,II31206,II31217,II31218,II31219,II31230,II31231,II31232,
    II31243,II31244,II31245,II31256,II31257,II31258,II31269,II31270,II31271,
    II31282,II31283,II31284,II31295,II31296,II31297,II31308,II31309,II31310,
    II31321,II31322,II31323,II31334,II31335,II31336,II31347,II31348,II31349,
    II31360,II31361,II31362,II31373,II31374,II31375,II31386,II31387,II31388,
    II31399,II31400,II31401,II31412,II31413,II31414,II31425,II31426,II31427,
    II31438,II31439,II31440,II31451,II31452,II31453,II31464,II31465,II31466,
    II31477,II31478,II31479,II31490,II31491,II31492,II31505,II31506,II31507,
    II31504,II31512,II31513,II31514,II31520,II31521,II31522,II31519,II31527,
    II31528,II31529,II31535,II31536,II31537,II31534,II31542,II31543,II31544,
    II31549,II31550,II31551,II31556,II31557,II31558,II31563,II31564,II31565,
    II31570,II31571,II31572,II31577,II31578,II31579,II31584,II31585,II31586,
    II31591,II31592,II31593,II31598,II31599,II31600,II31605,II31606,II31607,
    II31612,II31613,II31614,II31619,II31620,II31621,II31626,II31627,II31628,
    II31633,II31634,II31635,II31640,II31641,II31642,II31647,II31648,II31649,
    II31654,II31655,II31656,II31661,II31662,II31663,II31668,II31669,II31670,
    II31675,II31676,II31677,II31682,II31683,II31684,II31689,II31690,II31691,
    II31696,II31697,II31698,II31703,II31704,II31705,II31710,II31711,II31712,
    II31717,II31718,II31719,II31724,II31725,II31726,II31731,II31732,II31733,
    II31738,II31739,II31740,II31745,II31746,II31747,II34028,II34029,II34030,
    II34027,II34035,II34036,II34037,II34026,II34043,II34044,II34045,II34042,
    II34050,II34051,II34052,II34059,II34060,II34061,II34058,II34066,II34067,
    II34068,II34057,II34074,II34075,II34076,II34073,II34081,II34082,II34083,
    II34090,II34091,II34092,II34089,II34097,II34098,II34099,II34088,II34105,
    II34106,II34107,II34104,II34112,II34113,II34114,II34121,II34122,II34123,
    II34120,II34128,II34129,II34130,II34119,II34136,II34137,II34138,II34135,
    II34143,II34144,II34145,II34152,II34153,II34154,II34151,II34159,II34160,
    II34161,II34150,II34167,II34168,II34169,II34166,II34174,II34175,II34176,
    II34183,II34184,II34185,II34182,II34190,II34191,II34192,II34181,II34198,
    II34199,II34200,II34197,II34205,II34206,II34207,II34214,II34215,II34216,
    II34213,II34221,II34222,II34223,II34212,II34229,II34230,II34231,II34228,
    II34236,II34237,II34238,II34245,II34246,II34247,II34244,II34252,II34253,
    II34254,II34243,II34260,II34261,II34262,II34259,II34267,II34268,II34269,
    II34276,II34277,II34278,II34275,II34283,II34284,II34285,II34274,II34291,
    II34292,II34293,II34290,II34298,II34299,II34300,II34307,II34308,II34309,
    II34306,II34314,II34315,II34316,II34305,II34322,II34323,II34324,II34321,
    II34329,II34330,II34331,II34338,II34339,II34340,II34337,II34345,II34346,
    II34347,II34336,II34353,II34354,II34355,II34352,II34360,II34361,II34362,
    II34369,II34370,II34371,II34368,II34376,II34377,II34378,II34367,II34384,
    II34385,II34386,II34383,II34391,II34392,II34393,II34400,II34401,II34402,
    II34399,II34407,II34408,II34409,II34398,II34415,II34416,II34417,II34414,
    II34422,II34423,II34424,II34431,II34432,II34433,II34430,II34438,II34439,
    II34440,II34429,II34446,II34447,II34448,II34445,II34453,II34454,II34455,
    II34462,II34463,II34464,II34461,II34469,II34470,II34471,II34460,II34477,
    II34478,II34479,II34476,II34484,II34485,II34486,II34493,II34494,II34495,
    II34492,II34500,II34501,II34502,II34491,II34508,II34509,II34510,II34507,
    II34515,II34516,II34517,II34524,II34525,II34526,II34523,II34531,II34532,
    II34533,II34522,II34539,II34540,II34541,II34538,II34546,II34547,II34548,
    II34555,II34556,II34557,II34554,II34562,II34563,II34564,II34553,II34570,
    II34571,II34572,II34569,II34577,II34578,II34579,II34586,II34587,II34588,
    II34585,II34593,II34594,II34595,II34584,II34601,II34602,II34603,II34600,
    II34608,II34609,II34610,II34617,II34618,II34619,II34616,II34624,II34625,
    II34626,II34615,II34632,II34633,II34634,II34631,II34639,II34640,II34641,
    II34648,II34649,II34650,II34647,II34655,II34656,II34657,II34646,II34663,
    II34664,II34665,II34662,II34670,II34671,II34672,II34679,II34680,II34681,
    II34678,II34686,II34687,II34688,II34677,II34694,II34695,II34696,II34693,
    II34701,II34702,II34703,II34710,II34711,II34712,II34709,II34717,II34718,
    II34719,II34708,II34725,II34726,II34727,II34724,II34732,II34733,II34734,
    II34741,II34742,II34743,II34740,II34748,II34749,II34750,II34739,II34756,
    II34757,II34758,II34755,II34763,II34764,II34765,II34772,II34773,II34774,
    II34771,II34779,II34780,II34781,II34770,II34787,II34788,II34789,II34786,
    II34794,II34795,II34796,II34803,II34804,II34805,II34802,II34810,II34811,
    II34812,II34801,II34818,II34819,II34820,II34817,II34825,II34826,II34827,
    II34834,II34835,II34836,II34833,II34841,II34842,II34843,II34832,II34849,
    II34850,II34851,II34848,II34856,II34857,II34858,II34865,II34866,II34867,
    II34864,II34872,II34873,II34874,II34863,II34880,II34881,II34882,II34879,
    II34887,II34888,II34889,II34896,II34897,II34898,II34895,II34903,II34904,
    II34905,II34894,II34911,II34912,II34913,II34910,II34918,II34919,II34920,
    II34927,II34928,II34929,II34926,II34934,II34935,II34936,II34925,II34942,
    II34943,II34944,II34941,II34949,II34950,II34951,II34958,II34959,II34960,
    II34957,II34965,II34966,II34967,II34956,II34973,II34974,II34975,II34972,
    II34980,II34981,II34982,II34989,II34990,II34991,II34988,II34996,II34997,
    II34998,II34987,II35004,II35005,II35006,II35003,II35011,II35012,II35013,
    II35092,II35093,II35094,II35105,II35106,II35107,II35118,II35119,II35120,
    II35131,II35132,II35133,II35144,II35145,II35146,II35157,II35158,II35159,
    II35170,II35171,II35172,II35183,II35184,II35185,II35196,II35197,II35198,
    II35209,II35210,II35211,II35222,II35223,II35224,II35235,II35236,II35237,
    II35248,II35249,II35250,II35261,II35262,II35263,II35274,II35275,II35276,
    II35287,II35288,II35289,II35300,II35301,II35302,II35313,II35314,II35315,
    II35326,II35327,II35328,II35339,II35340,II35341,II35352,II35353,II35354,
    II35365,II35366,II35367,II35378,II35379,II35380,II35391,II35392,II35393,
    II35404,II35405,II35406,II35417,II35418,II35419,II35430,II35431,II35432,
    II35443,II35444,II35445,II35456,II35457,II35458,II35469,II35470,II35471,
    II35482,II35483,II35484,II35495,II35496,II35497,II35510,II35511,II35512,
    II35509,II35517,II35518,II35519,II35525,II35526,II35527,II35524,II35532,
    II35533,II35534,II35540,II35541,II35542,II35539,II35547,II35548,II35549,
    II35554,II35555,II35556,II35561,II35562,II35563,II35568,II35569,II35570,
    II35575,II35576,II35577,II35582,II35583,II35584,II35589,II35590,II35591,
    II35596,II35597,II35598,II35603,II35604,II35605,II35610,II35611,II35612,
    II35617,II35618,II35619,II35624,II35625,II35626,II35631,II35632,II35633,
    II35638,II35639,II35640,II35645,II35646,II35647,II35652,II35653,II35654,
    II35659,II35660,II35661,II35666,II35667,II35668,II35673,II35674,II35675,
    II35680,II35681,II35682,II35687,II35688,II35689,II35694,II35695,II35696,
    II35701,II35702,II35703,II35708,II35709,II35710,II35715,II35716,II35717,
    II35722,II35723,II35724,II35729,II35730,II35731,II35736,II35737,II35738,
    II35743,II35744,II35745,II35750,II35751,II35752;

  dff DFF_0(CK,WX485,WX484);
  dff DFF_1(CK,WX487,WX486);
  dff DFF_2(CK,WX489,WX488);
  dff DFF_3(CK,WX491,WX490);
  dff DFF_4(CK,WX493,WX492);
  dff DFF_5(CK,WX495,WX494);
  dff DFF_6(CK,WX497,WX496);
  dff DFF_7(CK,WX499,WX498);
  dff DFF_8(CK,WX501,WX500);
  dff DFF_9(CK,WX503,WX502);
  dff DFF_10(CK,WX505,WX504);
  dff DFF_11(CK,WX507,WX506);
  dff DFF_12(CK,WX509,WX508);
  dff DFF_13(CK,WX511,WX510);
  dff DFF_14(CK,WX513,WX512);
  dff DFF_15(CK,WX515,WX514);
  dff DFF_16(CK,WX517,WX516);
  dff DFF_17(CK,WX519,WX518);
  dff DFF_18(CK,WX521,WX520);
  dff DFF_19(CK,WX523,WX522);
  dff DFF_20(CK,WX525,WX524);
  dff DFF_21(CK,WX527,WX526);
  dff DFF_22(CK,WX529,WX528);
  dff DFF_23(CK,WX531,WX530);
  dff DFF_24(CK,WX533,WX532);
  dff DFF_25(CK,WX535,WX534);
  dff DFF_26(CK,WX537,WX536);
  dff DFF_27(CK,WX539,WX538);
  dff DFF_28(CK,WX541,WX540);
  dff DFF_29(CK,WX543,WX542);
  dff DFF_30(CK,WX545,WX544);
  dff DFF_31(CK,WX547,WX546);
  dff DFF_32(CK,WX645,WX644);
  dff DFF_33(CK,WX647,WX646);
  dff DFF_34(CK,WX649,WX648);
  dff DFF_35(CK,WX651,WX650);
  dff DFF_36(CK,WX653,WX652);
  dff DFF_37(CK,WX655,WX654);
  dff DFF_38(CK,WX657,WX656);
  dff DFF_39(CK,WX659,WX658);
  dff DFF_40(CK,WX661,WX660);
  dff DFF_41(CK,WX663,WX662);
  dff DFF_42(CK,WX665,WX664);
  dff DFF_43(CK,WX667,WX666);
  dff DFF_44(CK,WX669,WX668);
  dff DFF_45(CK,WX671,WX670);
  dff DFF_46(CK,WX673,WX672);
  dff DFF_47(CK,WX675,WX674);
  dff DFF_48(CK,WX677,WX676);
  dff DFF_49(CK,WX679,WX678);
  dff DFF_50(CK,WX681,WX680);
  dff DFF_51(CK,WX683,WX682);
  dff DFF_52(CK,WX685,WX684);
  dff DFF_53(CK,WX687,WX686);
  dff DFF_54(CK,WX689,WX688);
  dff DFF_55(CK,WX691,WX690);
  dff DFF_56(CK,WX693,WX692);
  dff DFF_57(CK,WX695,WX694);
  dff DFF_58(CK,WX697,WX696);
  dff DFF_59(CK,WX699,WX698);
  dff DFF_60(CK,WX701,WX700);
  dff DFF_61(CK,WX703,WX702);
  dff DFF_62(CK,WX705,WX704);
  dff DFF_63(CK,WX707,WX706);
  dff DFF_64(CK,WX709,WX708);
  dff DFF_65(CK,WX711,WX710);
  dff DFF_66(CK,WX713,WX712);
  dff DFF_67(CK,WX715,WX714);
  dff DFF_68(CK,WX717,WX716);
  dff DFF_69(CK,WX719,WX718);
  dff DFF_70(CK,WX721,WX720);
  dff DFF_71(CK,WX723,WX722);
  dff DFF_72(CK,WX725,WX724);
  dff DFF_73(CK,WX727,WX726);
  dff DFF_74(CK,WX729,WX728);
  dff DFF_75(CK,WX731,WX730);
  dff DFF_76(CK,WX733,WX732);
  dff DFF_77(CK,WX735,WX734);
  dff DFF_78(CK,WX737,WX736);
  dff DFF_79(CK,WX739,WX738);
  dff DFF_80(CK,WX741,WX740);
  dff DFF_81(CK,WX743,WX742);
  dff DFF_82(CK,WX745,WX744);
  dff DFF_83(CK,WX747,WX746);
  dff DFF_84(CK,WX749,WX748);
  dff DFF_85(CK,WX751,WX750);
  dff DFF_86(CK,WX753,WX752);
  dff DFF_87(CK,WX755,WX754);
  dff DFF_88(CK,WX757,WX756);
  dff DFF_89(CK,WX759,WX758);
  dff DFF_90(CK,WX761,WX760);
  dff DFF_91(CK,WX763,WX762);
  dff DFF_92(CK,WX765,WX764);
  dff DFF_93(CK,WX767,WX766);
  dff DFF_94(CK,WX769,WX768);
  dff DFF_95(CK,WX771,WX770);
  dff DFF_96(CK,WX773,WX772);
  dff DFF_97(CK,WX775,WX774);
  dff DFF_98(CK,WX777,WX776);
  dff DFF_99(CK,WX779,WX778);
  dff DFF_100(CK,WX781,WX780);
  dff DFF_101(CK,WX783,WX782);
  dff DFF_102(CK,WX785,WX784);
  dff DFF_103(CK,WX787,WX786);
  dff DFF_104(CK,WX789,WX788);
  dff DFF_105(CK,WX791,WX790);
  dff DFF_106(CK,WX793,WX792);
  dff DFF_107(CK,WX795,WX794);
  dff DFF_108(CK,WX797,WX796);
  dff DFF_109(CK,WX799,WX798);
  dff DFF_110(CK,WX801,WX800);
  dff DFF_111(CK,WX803,WX802);
  dff DFF_112(CK,WX805,WX804);
  dff DFF_113(CK,WX807,WX806);
  dff DFF_114(CK,WX809,WX808);
  dff DFF_115(CK,WX811,WX810);
  dff DFF_116(CK,WX813,WX812);
  dff DFF_117(CK,WX815,WX814);
  dff DFF_118(CK,WX817,WX816);
  dff DFF_119(CK,WX819,WX818);
  dff DFF_120(CK,WX821,WX820);
  dff DFF_121(CK,WX823,WX822);
  dff DFF_122(CK,WX825,WX824);
  dff DFF_123(CK,WX827,WX826);
  dff DFF_124(CK,WX829,WX828);
  dff DFF_125(CK,WX831,WX830);
  dff DFF_126(CK,WX833,WX832);
  dff DFF_127(CK,WX835,WX834);
  dff DFF_128(CK,WX837,WX836);
  dff DFF_129(CK,WX839,WX838);
  dff DFF_130(CK,WX841,WX840);
  dff DFF_131(CK,WX843,WX842);
  dff DFF_132(CK,WX845,WX844);
  dff DFF_133(CK,WX847,WX846);
  dff DFF_134(CK,WX849,WX848);
  dff DFF_135(CK,WX851,WX850);
  dff DFF_136(CK,WX853,WX852);
  dff DFF_137(CK,WX855,WX854);
  dff DFF_138(CK,WX857,WX856);
  dff DFF_139(CK,WX859,WX858);
  dff DFF_140(CK,WX861,WX860);
  dff DFF_141(CK,WX863,WX862);
  dff DFF_142(CK,WX865,WX864);
  dff DFF_143(CK,WX867,WX866);
  dff DFF_144(CK,WX869,WX868);
  dff DFF_145(CK,WX871,WX870);
  dff DFF_146(CK,WX873,WX872);
  dff DFF_147(CK,WX875,WX874);
  dff DFF_148(CK,WX877,WX876);
  dff DFF_149(CK,WX879,WX878);
  dff DFF_150(CK,WX881,WX880);
  dff DFF_151(CK,WX883,WX882);
  dff DFF_152(CK,WX885,WX884);
  dff DFF_153(CK,WX887,WX886);
  dff DFF_154(CK,WX889,WX888);
  dff DFF_155(CK,WX891,WX890);
  dff DFF_156(CK,WX893,WX892);
  dff DFF_157(CK,WX895,WX894);
  dff DFF_158(CK,WX897,WX896);
  dff DFF_159(CK,WX899,WX898);
  dff DFF_160(CK,CRC_OUT_9_0,WX1264);
  dff DFF_161(CK,CRC_OUT_9_1,WX1266);
  dff DFF_162(CK,CRC_OUT_9_2,WX1268);
  dff DFF_163(CK,CRC_OUT_9_3,WX1270);
  dff DFF_164(CK,CRC_OUT_9_4,WX1272);
  dff DFF_165(CK,CRC_OUT_9_5,WX1274);
  dff DFF_166(CK,CRC_OUT_9_6,WX1276);
  dff DFF_167(CK,CRC_OUT_9_7,WX1278);
  dff DFF_168(CK,CRC_OUT_9_8,WX1280);
  dff DFF_169(CK,CRC_OUT_9_9,WX1282);
  dff DFF_170(CK,CRC_OUT_9_10,WX1284);
  dff DFF_171(CK,CRC_OUT_9_11,WX1286);
  dff DFF_172(CK,CRC_OUT_9_12,WX1288);
  dff DFF_173(CK,CRC_OUT_9_13,WX1290);
  dff DFF_174(CK,CRC_OUT_9_14,WX1292);
  dff DFF_175(CK,CRC_OUT_9_15,WX1294);
  dff DFF_176(CK,CRC_OUT_9_16,WX1296);
  dff DFF_177(CK,CRC_OUT_9_17,WX1298);
  dff DFF_178(CK,CRC_OUT_9_18,WX1300);
  dff DFF_179(CK,CRC_OUT_9_19,WX1302);
  dff DFF_180(CK,CRC_OUT_9_20,WX1304);
  dff DFF_181(CK,CRC_OUT_9_21,WX1306);
  dff DFF_182(CK,CRC_OUT_9_22,WX1308);
  dff DFF_183(CK,CRC_OUT_9_23,WX1310);
  dff DFF_184(CK,CRC_OUT_9_24,WX1312);
  dff DFF_185(CK,CRC_OUT_9_25,WX1314);
  dff DFF_186(CK,CRC_OUT_9_26,WX1316);
  dff DFF_187(CK,CRC_OUT_9_27,WX1318);
  dff DFF_188(CK,CRC_OUT_9_28,WX1320);
  dff DFF_189(CK,CRC_OUT_9_29,WX1322);
  dff DFF_190(CK,CRC_OUT_9_30,WX1324);
  dff DFF_191(CK,CRC_OUT_9_31,WX1326);
  dff DFF_192(CK,WX1778,WX1777);
  dff DFF_193(CK,WX1780,WX1779);
  dff DFF_194(CK,WX1782,WX1781);
  dff DFF_195(CK,WX1784,WX1783);
  dff DFF_196(CK,WX1786,WX1785);
  dff DFF_197(CK,WX1788,WX1787);
  dff DFF_198(CK,WX1790,WX1789);
  dff DFF_199(CK,WX1792,WX1791);
  dff DFF_200(CK,WX1794,WX1793);
  dff DFF_201(CK,WX1796,WX1795);
  dff DFF_202(CK,WX1798,WX1797);
  dff DFF_203(CK,WX1800,WX1799);
  dff DFF_204(CK,WX1802,WX1801);
  dff DFF_205(CK,WX1804,WX1803);
  dff DFF_206(CK,WX1806,WX1805);
  dff DFF_207(CK,WX1808,WX1807);
  dff DFF_208(CK,WX1810,WX1809);
  dff DFF_209(CK,WX1812,WX1811);
  dff DFF_210(CK,WX1814,WX1813);
  dff DFF_211(CK,WX1816,WX1815);
  dff DFF_212(CK,WX1818,WX1817);
  dff DFF_213(CK,WX1820,WX1819);
  dff DFF_214(CK,WX1822,WX1821);
  dff DFF_215(CK,WX1824,WX1823);
  dff DFF_216(CK,WX1826,WX1825);
  dff DFF_217(CK,WX1828,WX1827);
  dff DFF_218(CK,WX1830,WX1829);
  dff DFF_219(CK,WX1832,WX1831);
  dff DFF_220(CK,WX1834,WX1833);
  dff DFF_221(CK,WX1836,WX1835);
  dff DFF_222(CK,WX1838,WX1837);
  dff DFF_223(CK,WX1840,WX1839);
  dff DFF_224(CK,WX1938,WX1937);
  dff DFF_225(CK,WX1940,WX1939);
  dff DFF_226(CK,WX1942,WX1941);
  dff DFF_227(CK,WX1944,WX1943);
  dff DFF_228(CK,WX1946,WX1945);
  dff DFF_229(CK,WX1948,WX1947);
  dff DFF_230(CK,WX1950,WX1949);
  dff DFF_231(CK,WX1952,WX1951);
  dff DFF_232(CK,WX1954,WX1953);
  dff DFF_233(CK,WX1956,WX1955);
  dff DFF_234(CK,WX1958,WX1957);
  dff DFF_235(CK,WX1960,WX1959);
  dff DFF_236(CK,WX1962,WX1961);
  dff DFF_237(CK,WX1964,WX1963);
  dff DFF_238(CK,WX1966,WX1965);
  dff DFF_239(CK,WX1968,WX1967);
  dff DFF_240(CK,WX1970,WX1969);
  dff DFF_241(CK,WX1972,WX1971);
  dff DFF_242(CK,WX1974,WX1973);
  dff DFF_243(CK,WX1976,WX1975);
  dff DFF_244(CK,WX1978,WX1977);
  dff DFF_245(CK,WX1980,WX1979);
  dff DFF_246(CK,WX1982,WX1981);
  dff DFF_247(CK,WX1984,WX1983);
  dff DFF_248(CK,WX1986,WX1985);
  dff DFF_249(CK,WX1988,WX1987);
  dff DFF_250(CK,WX1990,WX1989);
  dff DFF_251(CK,WX1992,WX1991);
  dff DFF_252(CK,WX1994,WX1993);
  dff DFF_253(CK,WX1996,WX1995);
  dff DFF_254(CK,WX1998,WX1997);
  dff DFF_255(CK,WX2000,WX1999);
  dff DFF_256(CK,WX2002,WX2001);
  dff DFF_257(CK,WX2004,WX2003);
  dff DFF_258(CK,WX2006,WX2005);
  dff DFF_259(CK,WX2008,WX2007);
  dff DFF_260(CK,WX2010,WX2009);
  dff DFF_261(CK,WX2012,WX2011);
  dff DFF_262(CK,WX2014,WX2013);
  dff DFF_263(CK,WX2016,WX2015);
  dff DFF_264(CK,WX2018,WX2017);
  dff DFF_265(CK,WX2020,WX2019);
  dff DFF_266(CK,WX2022,WX2021);
  dff DFF_267(CK,WX2024,WX2023);
  dff DFF_268(CK,WX2026,WX2025);
  dff DFF_269(CK,WX2028,WX2027);
  dff DFF_270(CK,WX2030,WX2029);
  dff DFF_271(CK,WX2032,WX2031);
  dff DFF_272(CK,WX2034,WX2033);
  dff DFF_273(CK,WX2036,WX2035);
  dff DFF_274(CK,WX2038,WX2037);
  dff DFF_275(CK,WX2040,WX2039);
  dff DFF_276(CK,WX2042,WX2041);
  dff DFF_277(CK,WX2044,WX2043);
  dff DFF_278(CK,WX2046,WX2045);
  dff DFF_279(CK,WX2048,WX2047);
  dff DFF_280(CK,WX2050,WX2049);
  dff DFF_281(CK,WX2052,WX2051);
  dff DFF_282(CK,WX2054,WX2053);
  dff DFF_283(CK,WX2056,WX2055);
  dff DFF_284(CK,WX2058,WX2057);
  dff DFF_285(CK,WX2060,WX2059);
  dff DFF_286(CK,WX2062,WX2061);
  dff DFF_287(CK,WX2064,WX2063);
  dff DFF_288(CK,WX2066,WX2065);
  dff DFF_289(CK,WX2068,WX2067);
  dff DFF_290(CK,WX2070,WX2069);
  dff DFF_291(CK,WX2072,WX2071);
  dff DFF_292(CK,WX2074,WX2073);
  dff DFF_293(CK,WX2076,WX2075);
  dff DFF_294(CK,WX2078,WX2077);
  dff DFF_295(CK,WX2080,WX2079);
  dff DFF_296(CK,WX2082,WX2081);
  dff DFF_297(CK,WX2084,WX2083);
  dff DFF_298(CK,WX2086,WX2085);
  dff DFF_299(CK,WX2088,WX2087);
  dff DFF_300(CK,WX2090,WX2089);
  dff DFF_301(CK,WX2092,WX2091);
  dff DFF_302(CK,WX2094,WX2093);
  dff DFF_303(CK,WX2096,WX2095);
  dff DFF_304(CK,WX2098,WX2097);
  dff DFF_305(CK,WX2100,WX2099);
  dff DFF_306(CK,WX2102,WX2101);
  dff DFF_307(CK,WX2104,WX2103);
  dff DFF_308(CK,WX2106,WX2105);
  dff DFF_309(CK,WX2108,WX2107);
  dff DFF_310(CK,WX2110,WX2109);
  dff DFF_311(CK,WX2112,WX2111);
  dff DFF_312(CK,WX2114,WX2113);
  dff DFF_313(CK,WX2116,WX2115);
  dff DFF_314(CK,WX2118,WX2117);
  dff DFF_315(CK,WX2120,WX2119);
  dff DFF_316(CK,WX2122,WX2121);
  dff DFF_317(CK,WX2124,WX2123);
  dff DFF_318(CK,WX2126,WX2125);
  dff DFF_319(CK,WX2128,WX2127);
  dff DFF_320(CK,WX2130,WX2129);
  dff DFF_321(CK,WX2132,WX2131);
  dff DFF_322(CK,WX2134,WX2133);
  dff DFF_323(CK,WX2136,WX2135);
  dff DFF_324(CK,WX2138,WX2137);
  dff DFF_325(CK,WX2140,WX2139);
  dff DFF_326(CK,WX2142,WX2141);
  dff DFF_327(CK,WX2144,WX2143);
  dff DFF_328(CK,WX2146,WX2145);
  dff DFF_329(CK,WX2148,WX2147);
  dff DFF_330(CK,WX2150,WX2149);
  dff DFF_331(CK,WX2152,WX2151);
  dff DFF_332(CK,WX2154,WX2153);
  dff DFF_333(CK,WX2156,WX2155);
  dff DFF_334(CK,WX2158,WX2157);
  dff DFF_335(CK,WX2160,WX2159);
  dff DFF_336(CK,WX2162,WX2161);
  dff DFF_337(CK,WX2164,WX2163);
  dff DFF_338(CK,WX2166,WX2165);
  dff DFF_339(CK,WX2168,WX2167);
  dff DFF_340(CK,WX2170,WX2169);
  dff DFF_341(CK,WX2172,WX2171);
  dff DFF_342(CK,WX2174,WX2173);
  dff DFF_343(CK,WX2176,WX2175);
  dff DFF_344(CK,WX2178,WX2177);
  dff DFF_345(CK,WX2180,WX2179);
  dff DFF_346(CK,WX2182,WX2181);
  dff DFF_347(CK,WX2184,WX2183);
  dff DFF_348(CK,WX2186,WX2185);
  dff DFF_349(CK,WX2188,WX2187);
  dff DFF_350(CK,WX2190,WX2189);
  dff DFF_351(CK,WX2192,WX2191);
  dff DFF_352(CK,CRC_OUT_8_0,WX2557);
  dff DFF_353(CK,CRC_OUT_8_1,WX2559);
  dff DFF_354(CK,CRC_OUT_8_2,WX2561);
  dff DFF_355(CK,CRC_OUT_8_3,WX2563);
  dff DFF_356(CK,CRC_OUT_8_4,WX2565);
  dff DFF_357(CK,CRC_OUT_8_5,WX2567);
  dff DFF_358(CK,CRC_OUT_8_6,WX2569);
  dff DFF_359(CK,CRC_OUT_8_7,WX2571);
  dff DFF_360(CK,CRC_OUT_8_8,WX2573);
  dff DFF_361(CK,CRC_OUT_8_9,WX2575);
  dff DFF_362(CK,CRC_OUT_8_10,WX2577);
  dff DFF_363(CK,CRC_OUT_8_11,WX2579);
  dff DFF_364(CK,CRC_OUT_8_12,WX2581);
  dff DFF_365(CK,CRC_OUT_8_13,WX2583);
  dff DFF_366(CK,CRC_OUT_8_14,WX2585);
  dff DFF_367(CK,CRC_OUT_8_15,WX2587);
  dff DFF_368(CK,CRC_OUT_8_16,WX2589);
  dff DFF_369(CK,CRC_OUT_8_17,WX2591);
  dff DFF_370(CK,CRC_OUT_8_18,WX2593);
  dff DFF_371(CK,CRC_OUT_8_19,WX2595);
  dff DFF_372(CK,CRC_OUT_8_20,WX2597);
  dff DFF_373(CK,CRC_OUT_8_21,WX2599);
  dff DFF_374(CK,CRC_OUT_8_22,WX2601);
  dff DFF_375(CK,CRC_OUT_8_23,WX2603);
  dff DFF_376(CK,CRC_OUT_8_24,WX2605);
  dff DFF_377(CK,CRC_OUT_8_25,WX2607);
  dff DFF_378(CK,CRC_OUT_8_26,WX2609);
  dff DFF_379(CK,CRC_OUT_8_27,WX2611);
  dff DFF_380(CK,CRC_OUT_8_28,WX2613);
  dff DFF_381(CK,CRC_OUT_8_29,WX2615);
  dff DFF_382(CK,CRC_OUT_8_30,WX2617);
  dff DFF_383(CK,CRC_OUT_8_31,WX2619);
  dff DFF_384(CK,WX3071,WX3070);
  dff DFF_385(CK,WX3073,WX3072);
  dff DFF_386(CK,WX3075,WX3074);
  dff DFF_387(CK,WX3077,WX3076);
  dff DFF_388(CK,WX3079,WX3078);
  dff DFF_389(CK,WX3081,WX3080);
  dff DFF_390(CK,WX3083,WX3082);
  dff DFF_391(CK,WX3085,WX3084);
  dff DFF_392(CK,WX3087,WX3086);
  dff DFF_393(CK,WX3089,WX3088);
  dff DFF_394(CK,WX3091,WX3090);
  dff DFF_395(CK,WX3093,WX3092);
  dff DFF_396(CK,WX3095,WX3094);
  dff DFF_397(CK,WX3097,WX3096);
  dff DFF_398(CK,WX3099,WX3098);
  dff DFF_399(CK,WX3101,WX3100);
  dff DFF_400(CK,WX3103,WX3102);
  dff DFF_401(CK,WX3105,WX3104);
  dff DFF_402(CK,WX3107,WX3106);
  dff DFF_403(CK,WX3109,WX3108);
  dff DFF_404(CK,WX3111,WX3110);
  dff DFF_405(CK,WX3113,WX3112);
  dff DFF_406(CK,WX3115,WX3114);
  dff DFF_407(CK,WX3117,WX3116);
  dff DFF_408(CK,WX3119,WX3118);
  dff DFF_409(CK,WX3121,WX3120);
  dff DFF_410(CK,WX3123,WX3122);
  dff DFF_411(CK,WX3125,WX3124);
  dff DFF_412(CK,WX3127,WX3126);
  dff DFF_413(CK,WX3129,WX3128);
  dff DFF_414(CK,WX3131,WX3130);
  dff DFF_415(CK,WX3133,WX3132);
  dff DFF_416(CK,WX3231,WX3230);
  dff DFF_417(CK,WX3233,WX3232);
  dff DFF_418(CK,WX3235,WX3234);
  dff DFF_419(CK,WX3237,WX3236);
  dff DFF_420(CK,WX3239,WX3238);
  dff DFF_421(CK,WX3241,WX3240);
  dff DFF_422(CK,WX3243,WX3242);
  dff DFF_423(CK,WX3245,WX3244);
  dff DFF_424(CK,WX3247,WX3246);
  dff DFF_425(CK,WX3249,WX3248);
  dff DFF_426(CK,WX3251,WX3250);
  dff DFF_427(CK,WX3253,WX3252);
  dff DFF_428(CK,WX3255,WX3254);
  dff DFF_429(CK,WX3257,WX3256);
  dff DFF_430(CK,WX3259,WX3258);
  dff DFF_431(CK,WX3261,WX3260);
  dff DFF_432(CK,WX3263,WX3262);
  dff DFF_433(CK,WX3265,WX3264);
  dff DFF_434(CK,WX3267,WX3266);
  dff DFF_435(CK,WX3269,WX3268);
  dff DFF_436(CK,WX3271,WX3270);
  dff DFF_437(CK,WX3273,WX3272);
  dff DFF_438(CK,WX3275,WX3274);
  dff DFF_439(CK,WX3277,WX3276);
  dff DFF_440(CK,WX3279,WX3278);
  dff DFF_441(CK,WX3281,WX3280);
  dff DFF_442(CK,WX3283,WX3282);
  dff DFF_443(CK,WX3285,WX3284);
  dff DFF_444(CK,WX3287,WX3286);
  dff DFF_445(CK,WX3289,WX3288);
  dff DFF_446(CK,WX3291,WX3290);
  dff DFF_447(CK,WX3293,WX3292);
  dff DFF_448(CK,WX3295,WX3294);
  dff DFF_449(CK,WX3297,WX3296);
  dff DFF_450(CK,WX3299,WX3298);
  dff DFF_451(CK,WX3301,WX3300);
  dff DFF_452(CK,WX3303,WX3302);
  dff DFF_453(CK,WX3305,WX3304);
  dff DFF_454(CK,WX3307,WX3306);
  dff DFF_455(CK,WX3309,WX3308);
  dff DFF_456(CK,WX3311,WX3310);
  dff DFF_457(CK,WX3313,WX3312);
  dff DFF_458(CK,WX3315,WX3314);
  dff DFF_459(CK,WX3317,WX3316);
  dff DFF_460(CK,WX3319,WX3318);
  dff DFF_461(CK,WX3321,WX3320);
  dff DFF_462(CK,WX3323,WX3322);
  dff DFF_463(CK,WX3325,WX3324);
  dff DFF_464(CK,WX3327,WX3326);
  dff DFF_465(CK,WX3329,WX3328);
  dff DFF_466(CK,WX3331,WX3330);
  dff DFF_467(CK,WX3333,WX3332);
  dff DFF_468(CK,WX3335,WX3334);
  dff DFF_469(CK,WX3337,WX3336);
  dff DFF_470(CK,WX3339,WX3338);
  dff DFF_471(CK,WX3341,WX3340);
  dff DFF_472(CK,WX3343,WX3342);
  dff DFF_473(CK,WX3345,WX3344);
  dff DFF_474(CK,WX3347,WX3346);
  dff DFF_475(CK,WX3349,WX3348);
  dff DFF_476(CK,WX3351,WX3350);
  dff DFF_477(CK,WX3353,WX3352);
  dff DFF_478(CK,WX3355,WX3354);
  dff DFF_479(CK,WX3357,WX3356);
  dff DFF_480(CK,WX3359,WX3358);
  dff DFF_481(CK,WX3361,WX3360);
  dff DFF_482(CK,WX3363,WX3362);
  dff DFF_483(CK,WX3365,WX3364);
  dff DFF_484(CK,WX3367,WX3366);
  dff DFF_485(CK,WX3369,WX3368);
  dff DFF_486(CK,WX3371,WX3370);
  dff DFF_487(CK,WX3373,WX3372);
  dff DFF_488(CK,WX3375,WX3374);
  dff DFF_489(CK,WX3377,WX3376);
  dff DFF_490(CK,WX3379,WX3378);
  dff DFF_491(CK,WX3381,WX3380);
  dff DFF_492(CK,WX3383,WX3382);
  dff DFF_493(CK,WX3385,WX3384);
  dff DFF_494(CK,WX3387,WX3386);
  dff DFF_495(CK,WX3389,WX3388);
  dff DFF_496(CK,WX3391,WX3390);
  dff DFF_497(CK,WX3393,WX3392);
  dff DFF_498(CK,WX3395,WX3394);
  dff DFF_499(CK,WX3397,WX3396);
  dff DFF_500(CK,WX3399,WX3398);
  dff DFF_501(CK,WX3401,WX3400);
  dff DFF_502(CK,WX3403,WX3402);
  dff DFF_503(CK,WX3405,WX3404);
  dff DFF_504(CK,WX3407,WX3406);
  dff DFF_505(CK,WX3409,WX3408);
  dff DFF_506(CK,WX3411,WX3410);
  dff DFF_507(CK,WX3413,WX3412);
  dff DFF_508(CK,WX3415,WX3414);
  dff DFF_509(CK,WX3417,WX3416);
  dff DFF_510(CK,WX3419,WX3418);
  dff DFF_511(CK,WX3421,WX3420);
  dff DFF_512(CK,WX3423,WX3422);
  dff DFF_513(CK,WX3425,WX3424);
  dff DFF_514(CK,WX3427,WX3426);
  dff DFF_515(CK,WX3429,WX3428);
  dff DFF_516(CK,WX3431,WX3430);
  dff DFF_517(CK,WX3433,WX3432);
  dff DFF_518(CK,WX3435,WX3434);
  dff DFF_519(CK,WX3437,WX3436);
  dff DFF_520(CK,WX3439,WX3438);
  dff DFF_521(CK,WX3441,WX3440);
  dff DFF_522(CK,WX3443,WX3442);
  dff DFF_523(CK,WX3445,WX3444);
  dff DFF_524(CK,WX3447,WX3446);
  dff DFF_525(CK,WX3449,WX3448);
  dff DFF_526(CK,WX3451,WX3450);
  dff DFF_527(CK,WX3453,WX3452);
  dff DFF_528(CK,WX3455,WX3454);
  dff DFF_529(CK,WX3457,WX3456);
  dff DFF_530(CK,WX3459,WX3458);
  dff DFF_531(CK,WX3461,WX3460);
  dff DFF_532(CK,WX3463,WX3462);
  dff DFF_533(CK,WX3465,WX3464);
  dff DFF_534(CK,WX3467,WX3466);
  dff DFF_535(CK,WX3469,WX3468);
  dff DFF_536(CK,WX3471,WX3470);
  dff DFF_537(CK,WX3473,WX3472);
  dff DFF_538(CK,WX3475,WX3474);
  dff DFF_539(CK,WX3477,WX3476);
  dff DFF_540(CK,WX3479,WX3478);
  dff DFF_541(CK,WX3481,WX3480);
  dff DFF_542(CK,WX3483,WX3482);
  dff DFF_543(CK,WX3485,WX3484);
  dff DFF_544(CK,CRC_OUT_7_0,WX3850);
  dff DFF_545(CK,CRC_OUT_7_1,WX3852);
  dff DFF_546(CK,CRC_OUT_7_2,WX3854);
  dff DFF_547(CK,CRC_OUT_7_3,WX3856);
  dff DFF_548(CK,CRC_OUT_7_4,WX3858);
  dff DFF_549(CK,CRC_OUT_7_5,WX3860);
  dff DFF_550(CK,CRC_OUT_7_6,WX3862);
  dff DFF_551(CK,CRC_OUT_7_7,WX3864);
  dff DFF_552(CK,CRC_OUT_7_8,WX3866);
  dff DFF_553(CK,CRC_OUT_7_9,WX3868);
  dff DFF_554(CK,CRC_OUT_7_10,WX3870);
  dff DFF_555(CK,CRC_OUT_7_11,WX3872);
  dff DFF_556(CK,CRC_OUT_7_12,WX3874);
  dff DFF_557(CK,CRC_OUT_7_13,WX3876);
  dff DFF_558(CK,CRC_OUT_7_14,WX3878);
  dff DFF_559(CK,CRC_OUT_7_15,WX3880);
  dff DFF_560(CK,CRC_OUT_7_16,WX3882);
  dff DFF_561(CK,CRC_OUT_7_17,WX3884);
  dff DFF_562(CK,CRC_OUT_7_18,WX3886);
  dff DFF_563(CK,CRC_OUT_7_19,WX3888);
  dff DFF_564(CK,CRC_OUT_7_20,WX3890);
  dff DFF_565(CK,CRC_OUT_7_21,WX3892);
  dff DFF_566(CK,CRC_OUT_7_22,WX3894);
  dff DFF_567(CK,CRC_OUT_7_23,WX3896);
  dff DFF_568(CK,CRC_OUT_7_24,WX3898);
  dff DFF_569(CK,CRC_OUT_7_25,WX3900);
  dff DFF_570(CK,CRC_OUT_7_26,WX3902);
  dff DFF_571(CK,CRC_OUT_7_27,WX3904);
  dff DFF_572(CK,CRC_OUT_7_28,WX3906);
  dff DFF_573(CK,CRC_OUT_7_29,WX3908);
  dff DFF_574(CK,CRC_OUT_7_30,WX3910);
  dff DFF_575(CK,CRC_OUT_7_31,WX3912);
  dff DFF_576(CK,WX4364,WX4363);
  dff DFF_577(CK,WX4366,WX4365);
  dff DFF_578(CK,WX4368,WX4367);
  dff DFF_579(CK,WX4370,WX4369);
  dff DFF_580(CK,WX4372,WX4371);
  dff DFF_581(CK,WX4374,WX4373);
  dff DFF_582(CK,WX4376,WX4375);
  dff DFF_583(CK,WX4378,WX4377);
  dff DFF_584(CK,WX4380,WX4379);
  dff DFF_585(CK,WX4382,WX4381);
  dff DFF_586(CK,WX4384,WX4383);
  dff DFF_587(CK,WX4386,WX4385);
  dff DFF_588(CK,WX4388,WX4387);
  dff DFF_589(CK,WX4390,WX4389);
  dff DFF_590(CK,WX4392,WX4391);
  dff DFF_591(CK,WX4394,WX4393);
  dff DFF_592(CK,WX4396,WX4395);
  dff DFF_593(CK,WX4398,WX4397);
  dff DFF_594(CK,WX4400,WX4399);
  dff DFF_595(CK,WX4402,WX4401);
  dff DFF_596(CK,WX4404,WX4403);
  dff DFF_597(CK,WX4406,WX4405);
  dff DFF_598(CK,WX4408,WX4407);
  dff DFF_599(CK,WX4410,WX4409);
  dff DFF_600(CK,WX4412,WX4411);
  dff DFF_601(CK,WX4414,WX4413);
  dff DFF_602(CK,WX4416,WX4415);
  dff DFF_603(CK,WX4418,WX4417);
  dff DFF_604(CK,WX4420,WX4419);
  dff DFF_605(CK,WX4422,WX4421);
  dff DFF_606(CK,WX4424,WX4423);
  dff DFF_607(CK,WX4426,WX4425);
  dff DFF_608(CK,WX4524,WX4523);
  dff DFF_609(CK,WX4526,WX4525);
  dff DFF_610(CK,WX4528,WX4527);
  dff DFF_611(CK,WX4530,WX4529);
  dff DFF_612(CK,WX4532,WX4531);
  dff DFF_613(CK,WX4534,WX4533);
  dff DFF_614(CK,WX4536,WX4535);
  dff DFF_615(CK,WX4538,WX4537);
  dff DFF_616(CK,WX4540,WX4539);
  dff DFF_617(CK,WX4542,WX4541);
  dff DFF_618(CK,WX4544,WX4543);
  dff DFF_619(CK,WX4546,WX4545);
  dff DFF_620(CK,WX4548,WX4547);
  dff DFF_621(CK,WX4550,WX4549);
  dff DFF_622(CK,WX4552,WX4551);
  dff DFF_623(CK,WX4554,WX4553);
  dff DFF_624(CK,WX4556,WX4555);
  dff DFF_625(CK,WX4558,WX4557);
  dff DFF_626(CK,WX4560,WX4559);
  dff DFF_627(CK,WX4562,WX4561);
  dff DFF_628(CK,WX4564,WX4563);
  dff DFF_629(CK,WX4566,WX4565);
  dff DFF_630(CK,WX4568,WX4567);
  dff DFF_631(CK,WX4570,WX4569);
  dff DFF_632(CK,WX4572,WX4571);
  dff DFF_633(CK,WX4574,WX4573);
  dff DFF_634(CK,WX4576,WX4575);
  dff DFF_635(CK,WX4578,WX4577);
  dff DFF_636(CK,WX4580,WX4579);
  dff DFF_637(CK,WX4582,WX4581);
  dff DFF_638(CK,WX4584,WX4583);
  dff DFF_639(CK,WX4586,WX4585);
  dff DFF_640(CK,WX4588,WX4587);
  dff DFF_641(CK,WX4590,WX4589);
  dff DFF_642(CK,WX4592,WX4591);
  dff DFF_643(CK,WX4594,WX4593);
  dff DFF_644(CK,WX4596,WX4595);
  dff DFF_645(CK,WX4598,WX4597);
  dff DFF_646(CK,WX4600,WX4599);
  dff DFF_647(CK,WX4602,WX4601);
  dff DFF_648(CK,WX4604,WX4603);
  dff DFF_649(CK,WX4606,WX4605);
  dff DFF_650(CK,WX4608,WX4607);
  dff DFF_651(CK,WX4610,WX4609);
  dff DFF_652(CK,WX4612,WX4611);
  dff DFF_653(CK,WX4614,WX4613);
  dff DFF_654(CK,WX4616,WX4615);
  dff DFF_655(CK,WX4618,WX4617);
  dff DFF_656(CK,WX4620,WX4619);
  dff DFF_657(CK,WX4622,WX4621);
  dff DFF_658(CK,WX4624,WX4623);
  dff DFF_659(CK,WX4626,WX4625);
  dff DFF_660(CK,WX4628,WX4627);
  dff DFF_661(CK,WX4630,WX4629);
  dff DFF_662(CK,WX4632,WX4631);
  dff DFF_663(CK,WX4634,WX4633);
  dff DFF_664(CK,WX4636,WX4635);
  dff DFF_665(CK,WX4638,WX4637);
  dff DFF_666(CK,WX4640,WX4639);
  dff DFF_667(CK,WX4642,WX4641);
  dff DFF_668(CK,WX4644,WX4643);
  dff DFF_669(CK,WX4646,WX4645);
  dff DFF_670(CK,WX4648,WX4647);
  dff DFF_671(CK,WX4650,WX4649);
  dff DFF_672(CK,WX4652,WX4651);
  dff DFF_673(CK,WX4654,WX4653);
  dff DFF_674(CK,WX4656,WX4655);
  dff DFF_675(CK,WX4658,WX4657);
  dff DFF_676(CK,WX4660,WX4659);
  dff DFF_677(CK,WX4662,WX4661);
  dff DFF_678(CK,WX4664,WX4663);
  dff DFF_679(CK,WX4666,WX4665);
  dff DFF_680(CK,WX4668,WX4667);
  dff DFF_681(CK,WX4670,WX4669);
  dff DFF_682(CK,WX4672,WX4671);
  dff DFF_683(CK,WX4674,WX4673);
  dff DFF_684(CK,WX4676,WX4675);
  dff DFF_685(CK,WX4678,WX4677);
  dff DFF_686(CK,WX4680,WX4679);
  dff DFF_687(CK,WX4682,WX4681);
  dff DFF_688(CK,WX4684,WX4683);
  dff DFF_689(CK,WX4686,WX4685);
  dff DFF_690(CK,WX4688,WX4687);
  dff DFF_691(CK,WX4690,WX4689);
  dff DFF_692(CK,WX4692,WX4691);
  dff DFF_693(CK,WX4694,WX4693);
  dff DFF_694(CK,WX4696,WX4695);
  dff DFF_695(CK,WX4698,WX4697);
  dff DFF_696(CK,WX4700,WX4699);
  dff DFF_697(CK,WX4702,WX4701);
  dff DFF_698(CK,WX4704,WX4703);
  dff DFF_699(CK,WX4706,WX4705);
  dff DFF_700(CK,WX4708,WX4707);
  dff DFF_701(CK,WX4710,WX4709);
  dff DFF_702(CK,WX4712,WX4711);
  dff DFF_703(CK,WX4714,WX4713);
  dff DFF_704(CK,WX4716,WX4715);
  dff DFF_705(CK,WX4718,WX4717);
  dff DFF_706(CK,WX4720,WX4719);
  dff DFF_707(CK,WX4722,WX4721);
  dff DFF_708(CK,WX4724,WX4723);
  dff DFF_709(CK,WX4726,WX4725);
  dff DFF_710(CK,WX4728,WX4727);
  dff DFF_711(CK,WX4730,WX4729);
  dff DFF_712(CK,WX4732,WX4731);
  dff DFF_713(CK,WX4734,WX4733);
  dff DFF_714(CK,WX4736,WX4735);
  dff DFF_715(CK,WX4738,WX4737);
  dff DFF_716(CK,WX4740,WX4739);
  dff DFF_717(CK,WX4742,WX4741);
  dff DFF_718(CK,WX4744,WX4743);
  dff DFF_719(CK,WX4746,WX4745);
  dff DFF_720(CK,WX4748,WX4747);
  dff DFF_721(CK,WX4750,WX4749);
  dff DFF_722(CK,WX4752,WX4751);
  dff DFF_723(CK,WX4754,WX4753);
  dff DFF_724(CK,WX4756,WX4755);
  dff DFF_725(CK,WX4758,WX4757);
  dff DFF_726(CK,WX4760,WX4759);
  dff DFF_727(CK,WX4762,WX4761);
  dff DFF_728(CK,WX4764,WX4763);
  dff DFF_729(CK,WX4766,WX4765);
  dff DFF_730(CK,WX4768,WX4767);
  dff DFF_731(CK,WX4770,WX4769);
  dff DFF_732(CK,WX4772,WX4771);
  dff DFF_733(CK,WX4774,WX4773);
  dff DFF_734(CK,WX4776,WX4775);
  dff DFF_735(CK,WX4778,WX4777);
  dff DFF_736(CK,CRC_OUT_6_0,WX5143);
  dff DFF_737(CK,CRC_OUT_6_1,WX5145);
  dff DFF_738(CK,CRC_OUT_6_2,WX5147);
  dff DFF_739(CK,CRC_OUT_6_3,WX5149);
  dff DFF_740(CK,CRC_OUT_6_4,WX5151);
  dff DFF_741(CK,CRC_OUT_6_5,WX5153);
  dff DFF_742(CK,CRC_OUT_6_6,WX5155);
  dff DFF_743(CK,CRC_OUT_6_7,WX5157);
  dff DFF_744(CK,CRC_OUT_6_8,WX5159);
  dff DFF_745(CK,CRC_OUT_6_9,WX5161);
  dff DFF_746(CK,CRC_OUT_6_10,WX5163);
  dff DFF_747(CK,CRC_OUT_6_11,WX5165);
  dff DFF_748(CK,CRC_OUT_6_12,WX5167);
  dff DFF_749(CK,CRC_OUT_6_13,WX5169);
  dff DFF_750(CK,CRC_OUT_6_14,WX5171);
  dff DFF_751(CK,CRC_OUT_6_15,WX5173);
  dff DFF_752(CK,CRC_OUT_6_16,WX5175);
  dff DFF_753(CK,CRC_OUT_6_17,WX5177);
  dff DFF_754(CK,CRC_OUT_6_18,WX5179);
  dff DFF_755(CK,CRC_OUT_6_19,WX5181);
  dff DFF_756(CK,CRC_OUT_6_20,WX5183);
  dff DFF_757(CK,CRC_OUT_6_21,WX5185);
  dff DFF_758(CK,CRC_OUT_6_22,WX5187);
  dff DFF_759(CK,CRC_OUT_6_23,WX5189);
  dff DFF_760(CK,CRC_OUT_6_24,WX5191);
  dff DFF_761(CK,CRC_OUT_6_25,WX5193);
  dff DFF_762(CK,CRC_OUT_6_26,WX5195);
  dff DFF_763(CK,CRC_OUT_6_27,WX5197);
  dff DFF_764(CK,CRC_OUT_6_28,WX5199);
  dff DFF_765(CK,CRC_OUT_6_29,WX5201);
  dff DFF_766(CK,CRC_OUT_6_30,WX5203);
  dff DFF_767(CK,CRC_OUT_6_31,WX5205);
  dff DFF_768(CK,WX5657,WX5656);
  dff DFF_769(CK,WX5659,WX5658);
  dff DFF_770(CK,WX5661,WX5660);
  dff DFF_771(CK,WX5663,WX5662);
  dff DFF_772(CK,WX5665,WX5664);
  dff DFF_773(CK,WX5667,WX5666);
  dff DFF_774(CK,WX5669,WX5668);
  dff DFF_775(CK,WX5671,WX5670);
  dff DFF_776(CK,WX5673,WX5672);
  dff DFF_777(CK,WX5675,WX5674);
  dff DFF_778(CK,WX5677,WX5676);
  dff DFF_779(CK,WX5679,WX5678);
  dff DFF_780(CK,WX5681,WX5680);
  dff DFF_781(CK,WX5683,WX5682);
  dff DFF_782(CK,WX5685,WX5684);
  dff DFF_783(CK,WX5687,WX5686);
  dff DFF_784(CK,WX5689,WX5688);
  dff DFF_785(CK,WX5691,WX5690);
  dff DFF_786(CK,WX5693,WX5692);
  dff DFF_787(CK,WX5695,WX5694);
  dff DFF_788(CK,WX5697,WX5696);
  dff DFF_789(CK,WX5699,WX5698);
  dff DFF_790(CK,WX5701,WX5700);
  dff DFF_791(CK,WX5703,WX5702);
  dff DFF_792(CK,WX5705,WX5704);
  dff DFF_793(CK,WX5707,WX5706);
  dff DFF_794(CK,WX5709,WX5708);
  dff DFF_795(CK,WX5711,WX5710);
  dff DFF_796(CK,WX5713,WX5712);
  dff DFF_797(CK,WX5715,WX5714);
  dff DFF_798(CK,WX5717,WX5716);
  dff DFF_799(CK,WX5719,WX5718);
  dff DFF_800(CK,WX5817,WX5816);
  dff DFF_801(CK,WX5819,WX5818);
  dff DFF_802(CK,WX5821,WX5820);
  dff DFF_803(CK,WX5823,WX5822);
  dff DFF_804(CK,WX5825,WX5824);
  dff DFF_805(CK,WX5827,WX5826);
  dff DFF_806(CK,WX5829,WX5828);
  dff DFF_807(CK,WX5831,WX5830);
  dff DFF_808(CK,WX5833,WX5832);
  dff DFF_809(CK,WX5835,WX5834);
  dff DFF_810(CK,WX5837,WX5836);
  dff DFF_811(CK,WX5839,WX5838);
  dff DFF_812(CK,WX5841,WX5840);
  dff DFF_813(CK,WX5843,WX5842);
  dff DFF_814(CK,WX5845,WX5844);
  dff DFF_815(CK,WX5847,WX5846);
  dff DFF_816(CK,WX5849,WX5848);
  dff DFF_817(CK,WX5851,WX5850);
  dff DFF_818(CK,WX5853,WX5852);
  dff DFF_819(CK,WX5855,WX5854);
  dff DFF_820(CK,WX5857,WX5856);
  dff DFF_821(CK,WX5859,WX5858);
  dff DFF_822(CK,WX5861,WX5860);
  dff DFF_823(CK,WX5863,WX5862);
  dff DFF_824(CK,WX5865,WX5864);
  dff DFF_825(CK,WX5867,WX5866);
  dff DFF_826(CK,WX5869,WX5868);
  dff DFF_827(CK,WX5871,WX5870);
  dff DFF_828(CK,WX5873,WX5872);
  dff DFF_829(CK,WX5875,WX5874);
  dff DFF_830(CK,WX5877,WX5876);
  dff DFF_831(CK,WX5879,WX5878);
  dff DFF_832(CK,WX5881,WX5880);
  dff DFF_833(CK,WX5883,WX5882);
  dff DFF_834(CK,WX5885,WX5884);
  dff DFF_835(CK,WX5887,WX5886);
  dff DFF_836(CK,WX5889,WX5888);
  dff DFF_837(CK,WX5891,WX5890);
  dff DFF_838(CK,WX5893,WX5892);
  dff DFF_839(CK,WX5895,WX5894);
  dff DFF_840(CK,WX5897,WX5896);
  dff DFF_841(CK,WX5899,WX5898);
  dff DFF_842(CK,WX5901,WX5900);
  dff DFF_843(CK,WX5903,WX5902);
  dff DFF_844(CK,WX5905,WX5904);
  dff DFF_845(CK,WX5907,WX5906);
  dff DFF_846(CK,WX5909,WX5908);
  dff DFF_847(CK,WX5911,WX5910);
  dff DFF_848(CK,WX5913,WX5912);
  dff DFF_849(CK,WX5915,WX5914);
  dff DFF_850(CK,WX5917,WX5916);
  dff DFF_851(CK,WX5919,WX5918);
  dff DFF_852(CK,WX5921,WX5920);
  dff DFF_853(CK,WX5923,WX5922);
  dff DFF_854(CK,WX5925,WX5924);
  dff DFF_855(CK,WX5927,WX5926);
  dff DFF_856(CK,WX5929,WX5928);
  dff DFF_857(CK,WX5931,WX5930);
  dff DFF_858(CK,WX5933,WX5932);
  dff DFF_859(CK,WX5935,WX5934);
  dff DFF_860(CK,WX5937,WX5936);
  dff DFF_861(CK,WX5939,WX5938);
  dff DFF_862(CK,WX5941,WX5940);
  dff DFF_863(CK,WX5943,WX5942);
  dff DFF_864(CK,WX5945,WX5944);
  dff DFF_865(CK,WX5947,WX5946);
  dff DFF_866(CK,WX5949,WX5948);
  dff DFF_867(CK,WX5951,WX5950);
  dff DFF_868(CK,WX5953,WX5952);
  dff DFF_869(CK,WX5955,WX5954);
  dff DFF_870(CK,WX5957,WX5956);
  dff DFF_871(CK,WX5959,WX5958);
  dff DFF_872(CK,WX5961,WX5960);
  dff DFF_873(CK,WX5963,WX5962);
  dff DFF_874(CK,WX5965,WX5964);
  dff DFF_875(CK,WX5967,WX5966);
  dff DFF_876(CK,WX5969,WX5968);
  dff DFF_877(CK,WX5971,WX5970);
  dff DFF_878(CK,WX5973,WX5972);
  dff DFF_879(CK,WX5975,WX5974);
  dff DFF_880(CK,WX5977,WX5976);
  dff DFF_881(CK,WX5979,WX5978);
  dff DFF_882(CK,WX5981,WX5980);
  dff DFF_883(CK,WX5983,WX5982);
  dff DFF_884(CK,WX5985,WX5984);
  dff DFF_885(CK,WX5987,WX5986);
  dff DFF_886(CK,WX5989,WX5988);
  dff DFF_887(CK,WX5991,WX5990);
  dff DFF_888(CK,WX5993,WX5992);
  dff DFF_889(CK,WX5995,WX5994);
  dff DFF_890(CK,WX5997,WX5996);
  dff DFF_891(CK,WX5999,WX5998);
  dff DFF_892(CK,WX6001,WX6000);
  dff DFF_893(CK,WX6003,WX6002);
  dff DFF_894(CK,WX6005,WX6004);
  dff DFF_895(CK,WX6007,WX6006);
  dff DFF_896(CK,WX6009,WX6008);
  dff DFF_897(CK,WX6011,WX6010);
  dff DFF_898(CK,WX6013,WX6012);
  dff DFF_899(CK,WX6015,WX6014);
  dff DFF_900(CK,WX6017,WX6016);
  dff DFF_901(CK,WX6019,WX6018);
  dff DFF_902(CK,WX6021,WX6020);
  dff DFF_903(CK,WX6023,WX6022);
  dff DFF_904(CK,WX6025,WX6024);
  dff DFF_905(CK,WX6027,WX6026);
  dff DFF_906(CK,WX6029,WX6028);
  dff DFF_907(CK,WX6031,WX6030);
  dff DFF_908(CK,WX6033,WX6032);
  dff DFF_909(CK,WX6035,WX6034);
  dff DFF_910(CK,WX6037,WX6036);
  dff DFF_911(CK,WX6039,WX6038);
  dff DFF_912(CK,WX6041,WX6040);
  dff DFF_913(CK,WX6043,WX6042);
  dff DFF_914(CK,WX6045,WX6044);
  dff DFF_915(CK,WX6047,WX6046);
  dff DFF_916(CK,WX6049,WX6048);
  dff DFF_917(CK,WX6051,WX6050);
  dff DFF_918(CK,WX6053,WX6052);
  dff DFF_919(CK,WX6055,WX6054);
  dff DFF_920(CK,WX6057,WX6056);
  dff DFF_921(CK,WX6059,WX6058);
  dff DFF_922(CK,WX6061,WX6060);
  dff DFF_923(CK,WX6063,WX6062);
  dff DFF_924(CK,WX6065,WX6064);
  dff DFF_925(CK,WX6067,WX6066);
  dff DFF_926(CK,WX6069,WX6068);
  dff DFF_927(CK,WX6071,WX6070);
  dff DFF_928(CK,CRC_OUT_5_0,WX6436);
  dff DFF_929(CK,CRC_OUT_5_1,WX6438);
  dff DFF_930(CK,CRC_OUT_5_2,WX6440);
  dff DFF_931(CK,CRC_OUT_5_3,WX6442);
  dff DFF_932(CK,CRC_OUT_5_4,WX6444);
  dff DFF_933(CK,CRC_OUT_5_5,WX6446);
  dff DFF_934(CK,CRC_OUT_5_6,WX6448);
  dff DFF_935(CK,CRC_OUT_5_7,WX6450);
  dff DFF_936(CK,CRC_OUT_5_8,WX6452);
  dff DFF_937(CK,CRC_OUT_5_9,WX6454);
  dff DFF_938(CK,CRC_OUT_5_10,WX6456);
  dff DFF_939(CK,CRC_OUT_5_11,WX6458);
  dff DFF_940(CK,CRC_OUT_5_12,WX6460);
  dff DFF_941(CK,CRC_OUT_5_13,WX6462);
  dff DFF_942(CK,CRC_OUT_5_14,WX6464);
  dff DFF_943(CK,CRC_OUT_5_15,WX6466);
  dff DFF_944(CK,CRC_OUT_5_16,WX6468);
  dff DFF_945(CK,CRC_OUT_5_17,WX6470);
  dff DFF_946(CK,CRC_OUT_5_18,WX6472);
  dff DFF_947(CK,CRC_OUT_5_19,WX6474);
  dff DFF_948(CK,CRC_OUT_5_20,WX6476);
  dff DFF_949(CK,CRC_OUT_5_21,WX6478);
  dff DFF_950(CK,CRC_OUT_5_22,WX6480);
  dff DFF_951(CK,CRC_OUT_5_23,WX6482);
  dff DFF_952(CK,CRC_OUT_5_24,WX6484);
  dff DFF_953(CK,CRC_OUT_5_25,WX6486);
  dff DFF_954(CK,CRC_OUT_5_26,WX6488);
  dff DFF_955(CK,CRC_OUT_5_27,WX6490);
  dff DFF_956(CK,CRC_OUT_5_28,WX6492);
  dff DFF_957(CK,CRC_OUT_5_29,WX6494);
  dff DFF_958(CK,CRC_OUT_5_30,WX6496);
  dff DFF_959(CK,CRC_OUT_5_31,WX6498);
  dff DFF_960(CK,WX6950,WX6949);
  dff DFF_961(CK,WX6952,WX6951);
  dff DFF_962(CK,WX6954,WX6953);
  dff DFF_963(CK,WX6956,WX6955);
  dff DFF_964(CK,WX6958,WX6957);
  dff DFF_965(CK,WX6960,WX6959);
  dff DFF_966(CK,WX6962,WX6961);
  dff DFF_967(CK,WX6964,WX6963);
  dff DFF_968(CK,WX6966,WX6965);
  dff DFF_969(CK,WX6968,WX6967);
  dff DFF_970(CK,WX6970,WX6969);
  dff DFF_971(CK,WX6972,WX6971);
  dff DFF_972(CK,WX6974,WX6973);
  dff DFF_973(CK,WX6976,WX6975);
  dff DFF_974(CK,WX6978,WX6977);
  dff DFF_975(CK,WX6980,WX6979);
  dff DFF_976(CK,WX6982,WX6981);
  dff DFF_977(CK,WX6984,WX6983);
  dff DFF_978(CK,WX6986,WX6985);
  dff DFF_979(CK,WX6988,WX6987);
  dff DFF_980(CK,WX6990,WX6989);
  dff DFF_981(CK,WX6992,WX6991);
  dff DFF_982(CK,WX6994,WX6993);
  dff DFF_983(CK,WX6996,WX6995);
  dff DFF_984(CK,WX6998,WX6997);
  dff DFF_985(CK,WX7000,WX6999);
  dff DFF_986(CK,WX7002,WX7001);
  dff DFF_987(CK,WX7004,WX7003);
  dff DFF_988(CK,WX7006,WX7005);
  dff DFF_989(CK,WX7008,WX7007);
  dff DFF_990(CK,WX7010,WX7009);
  dff DFF_991(CK,WX7012,WX7011);
  dff DFF_992(CK,WX7110,WX7109);
  dff DFF_993(CK,WX7112,WX7111);
  dff DFF_994(CK,WX7114,WX7113);
  dff DFF_995(CK,WX7116,WX7115);
  dff DFF_996(CK,WX7118,WX7117);
  dff DFF_997(CK,WX7120,WX7119);
  dff DFF_998(CK,WX7122,WX7121);
  dff DFF_999(CK,WX7124,WX7123);
  dff DFF_1000(CK,WX7126,WX7125);
  dff DFF_1001(CK,WX7128,WX7127);
  dff DFF_1002(CK,WX7130,WX7129);
  dff DFF_1003(CK,WX7132,WX7131);
  dff DFF_1004(CK,WX7134,WX7133);
  dff DFF_1005(CK,WX7136,WX7135);
  dff DFF_1006(CK,WX7138,WX7137);
  dff DFF_1007(CK,WX7140,WX7139);
  dff DFF_1008(CK,WX7142,WX7141);
  dff DFF_1009(CK,WX7144,WX7143);
  dff DFF_1010(CK,WX7146,WX7145);
  dff DFF_1011(CK,WX7148,WX7147);
  dff DFF_1012(CK,WX7150,WX7149);
  dff DFF_1013(CK,WX7152,WX7151);
  dff DFF_1014(CK,WX7154,WX7153);
  dff DFF_1015(CK,WX7156,WX7155);
  dff DFF_1016(CK,WX7158,WX7157);
  dff DFF_1017(CK,WX7160,WX7159);
  dff DFF_1018(CK,WX7162,WX7161);
  dff DFF_1019(CK,WX7164,WX7163);
  dff DFF_1020(CK,WX7166,WX7165);
  dff DFF_1021(CK,WX7168,WX7167);
  dff DFF_1022(CK,WX7170,WX7169);
  dff DFF_1023(CK,WX7172,WX7171);
  dff DFF_1024(CK,WX7174,WX7173);
  dff DFF_1025(CK,WX7176,WX7175);
  dff DFF_1026(CK,WX7178,WX7177);
  dff DFF_1027(CK,WX7180,WX7179);
  dff DFF_1028(CK,WX7182,WX7181);
  dff DFF_1029(CK,WX7184,WX7183);
  dff DFF_1030(CK,WX7186,WX7185);
  dff DFF_1031(CK,WX7188,WX7187);
  dff DFF_1032(CK,WX7190,WX7189);
  dff DFF_1033(CK,WX7192,WX7191);
  dff DFF_1034(CK,WX7194,WX7193);
  dff DFF_1035(CK,WX7196,WX7195);
  dff DFF_1036(CK,WX7198,WX7197);
  dff DFF_1037(CK,WX7200,WX7199);
  dff DFF_1038(CK,WX7202,WX7201);
  dff DFF_1039(CK,WX7204,WX7203);
  dff DFF_1040(CK,WX7206,WX7205);
  dff DFF_1041(CK,WX7208,WX7207);
  dff DFF_1042(CK,WX7210,WX7209);
  dff DFF_1043(CK,WX7212,WX7211);
  dff DFF_1044(CK,WX7214,WX7213);
  dff DFF_1045(CK,WX7216,WX7215);
  dff DFF_1046(CK,WX7218,WX7217);
  dff DFF_1047(CK,WX7220,WX7219);
  dff DFF_1048(CK,WX7222,WX7221);
  dff DFF_1049(CK,WX7224,WX7223);
  dff DFF_1050(CK,WX7226,WX7225);
  dff DFF_1051(CK,WX7228,WX7227);
  dff DFF_1052(CK,WX7230,WX7229);
  dff DFF_1053(CK,WX7232,WX7231);
  dff DFF_1054(CK,WX7234,WX7233);
  dff DFF_1055(CK,WX7236,WX7235);
  dff DFF_1056(CK,WX7238,WX7237);
  dff DFF_1057(CK,WX7240,WX7239);
  dff DFF_1058(CK,WX7242,WX7241);
  dff DFF_1059(CK,WX7244,WX7243);
  dff DFF_1060(CK,WX7246,WX7245);
  dff DFF_1061(CK,WX7248,WX7247);
  dff DFF_1062(CK,WX7250,WX7249);
  dff DFF_1063(CK,WX7252,WX7251);
  dff DFF_1064(CK,WX7254,WX7253);
  dff DFF_1065(CK,WX7256,WX7255);
  dff DFF_1066(CK,WX7258,WX7257);
  dff DFF_1067(CK,WX7260,WX7259);
  dff DFF_1068(CK,WX7262,WX7261);
  dff DFF_1069(CK,WX7264,WX7263);
  dff DFF_1070(CK,WX7266,WX7265);
  dff DFF_1071(CK,WX7268,WX7267);
  dff DFF_1072(CK,WX7270,WX7269);
  dff DFF_1073(CK,WX7272,WX7271);
  dff DFF_1074(CK,WX7274,WX7273);
  dff DFF_1075(CK,WX7276,WX7275);
  dff DFF_1076(CK,WX7278,WX7277);
  dff DFF_1077(CK,WX7280,WX7279);
  dff DFF_1078(CK,WX7282,WX7281);
  dff DFF_1079(CK,WX7284,WX7283);
  dff DFF_1080(CK,WX7286,WX7285);
  dff DFF_1081(CK,WX7288,WX7287);
  dff DFF_1082(CK,WX7290,WX7289);
  dff DFF_1083(CK,WX7292,WX7291);
  dff DFF_1084(CK,WX7294,WX7293);
  dff DFF_1085(CK,WX7296,WX7295);
  dff DFF_1086(CK,WX7298,WX7297);
  dff DFF_1087(CK,WX7300,WX7299);
  dff DFF_1088(CK,WX7302,WX7301);
  dff DFF_1089(CK,WX7304,WX7303);
  dff DFF_1090(CK,WX7306,WX7305);
  dff DFF_1091(CK,WX7308,WX7307);
  dff DFF_1092(CK,WX7310,WX7309);
  dff DFF_1093(CK,WX7312,WX7311);
  dff DFF_1094(CK,WX7314,WX7313);
  dff DFF_1095(CK,WX7316,WX7315);
  dff DFF_1096(CK,WX7318,WX7317);
  dff DFF_1097(CK,WX7320,WX7319);
  dff DFF_1098(CK,WX7322,WX7321);
  dff DFF_1099(CK,WX7324,WX7323);
  dff DFF_1100(CK,WX7326,WX7325);
  dff DFF_1101(CK,WX7328,WX7327);
  dff DFF_1102(CK,WX7330,WX7329);
  dff DFF_1103(CK,WX7332,WX7331);
  dff DFF_1104(CK,WX7334,WX7333);
  dff DFF_1105(CK,WX7336,WX7335);
  dff DFF_1106(CK,WX7338,WX7337);
  dff DFF_1107(CK,WX7340,WX7339);
  dff DFF_1108(CK,WX7342,WX7341);
  dff DFF_1109(CK,WX7344,WX7343);
  dff DFF_1110(CK,WX7346,WX7345);
  dff DFF_1111(CK,WX7348,WX7347);
  dff DFF_1112(CK,WX7350,WX7349);
  dff DFF_1113(CK,WX7352,WX7351);
  dff DFF_1114(CK,WX7354,WX7353);
  dff DFF_1115(CK,WX7356,WX7355);
  dff DFF_1116(CK,WX7358,WX7357);
  dff DFF_1117(CK,WX7360,WX7359);
  dff DFF_1118(CK,WX7362,WX7361);
  dff DFF_1119(CK,WX7364,WX7363);
  dff DFF_1120(CK,CRC_OUT_4_0,WX7729);
  dff DFF_1121(CK,CRC_OUT_4_1,WX7731);
  dff DFF_1122(CK,CRC_OUT_4_2,WX7733);
  dff DFF_1123(CK,CRC_OUT_4_3,WX7735);
  dff DFF_1124(CK,CRC_OUT_4_4,WX7737);
  dff DFF_1125(CK,CRC_OUT_4_5,WX7739);
  dff DFF_1126(CK,CRC_OUT_4_6,WX7741);
  dff DFF_1127(CK,CRC_OUT_4_7,WX7743);
  dff DFF_1128(CK,CRC_OUT_4_8,WX7745);
  dff DFF_1129(CK,CRC_OUT_4_9,WX7747);
  dff DFF_1130(CK,CRC_OUT_4_10,WX7749);
  dff DFF_1131(CK,CRC_OUT_4_11,WX7751);
  dff DFF_1132(CK,CRC_OUT_4_12,WX7753);
  dff DFF_1133(CK,CRC_OUT_4_13,WX7755);
  dff DFF_1134(CK,CRC_OUT_4_14,WX7757);
  dff DFF_1135(CK,CRC_OUT_4_15,WX7759);
  dff DFF_1136(CK,CRC_OUT_4_16,WX7761);
  dff DFF_1137(CK,CRC_OUT_4_17,WX7763);
  dff DFF_1138(CK,CRC_OUT_4_18,WX7765);
  dff DFF_1139(CK,CRC_OUT_4_19,WX7767);
  dff DFF_1140(CK,CRC_OUT_4_20,WX7769);
  dff DFF_1141(CK,CRC_OUT_4_21,WX7771);
  dff DFF_1142(CK,CRC_OUT_4_22,WX7773);
  dff DFF_1143(CK,CRC_OUT_4_23,WX7775);
  dff DFF_1144(CK,CRC_OUT_4_24,WX7777);
  dff DFF_1145(CK,CRC_OUT_4_25,WX7779);
  dff DFF_1146(CK,CRC_OUT_4_26,WX7781);
  dff DFF_1147(CK,CRC_OUT_4_27,WX7783);
  dff DFF_1148(CK,CRC_OUT_4_28,WX7785);
  dff DFF_1149(CK,CRC_OUT_4_29,WX7787);
  dff DFF_1150(CK,CRC_OUT_4_30,WX7789);
  dff DFF_1151(CK,CRC_OUT_4_31,WX7791);
  dff DFF_1152(CK,WX8243,WX8242);
  dff DFF_1153(CK,WX8245,WX8244);
  dff DFF_1154(CK,WX8247,WX8246);
  dff DFF_1155(CK,WX8249,WX8248);
  dff DFF_1156(CK,WX8251,WX8250);
  dff DFF_1157(CK,WX8253,WX8252);
  dff DFF_1158(CK,WX8255,WX8254);
  dff DFF_1159(CK,WX8257,WX8256);
  dff DFF_1160(CK,WX8259,WX8258);
  dff DFF_1161(CK,WX8261,WX8260);
  dff DFF_1162(CK,WX8263,WX8262);
  dff DFF_1163(CK,WX8265,WX8264);
  dff DFF_1164(CK,WX8267,WX8266);
  dff DFF_1165(CK,WX8269,WX8268);
  dff DFF_1166(CK,WX8271,WX8270);
  dff DFF_1167(CK,WX8273,WX8272);
  dff DFF_1168(CK,WX8275,WX8274);
  dff DFF_1169(CK,WX8277,WX8276);
  dff DFF_1170(CK,WX8279,WX8278);
  dff DFF_1171(CK,WX8281,WX8280);
  dff DFF_1172(CK,WX8283,WX8282);
  dff DFF_1173(CK,WX8285,WX8284);
  dff DFF_1174(CK,WX8287,WX8286);
  dff DFF_1175(CK,WX8289,WX8288);
  dff DFF_1176(CK,WX8291,WX8290);
  dff DFF_1177(CK,WX8293,WX8292);
  dff DFF_1178(CK,WX8295,WX8294);
  dff DFF_1179(CK,WX8297,WX8296);
  dff DFF_1180(CK,WX8299,WX8298);
  dff DFF_1181(CK,WX8301,WX8300);
  dff DFF_1182(CK,WX8303,WX8302);
  dff DFF_1183(CK,WX8305,WX8304);
  dff DFF_1184(CK,WX8403,WX8402);
  dff DFF_1185(CK,WX8405,WX8404);
  dff DFF_1186(CK,WX8407,WX8406);
  dff DFF_1187(CK,WX8409,WX8408);
  dff DFF_1188(CK,WX8411,WX8410);
  dff DFF_1189(CK,WX8413,WX8412);
  dff DFF_1190(CK,WX8415,WX8414);
  dff DFF_1191(CK,WX8417,WX8416);
  dff DFF_1192(CK,WX8419,WX8418);
  dff DFF_1193(CK,WX8421,WX8420);
  dff DFF_1194(CK,WX8423,WX8422);
  dff DFF_1195(CK,WX8425,WX8424);
  dff DFF_1196(CK,WX8427,WX8426);
  dff DFF_1197(CK,WX8429,WX8428);
  dff DFF_1198(CK,WX8431,WX8430);
  dff DFF_1199(CK,WX8433,WX8432);
  dff DFF_1200(CK,WX8435,WX8434);
  dff DFF_1201(CK,WX8437,WX8436);
  dff DFF_1202(CK,WX8439,WX8438);
  dff DFF_1203(CK,WX8441,WX8440);
  dff DFF_1204(CK,WX8443,WX8442);
  dff DFF_1205(CK,WX8445,WX8444);
  dff DFF_1206(CK,WX8447,WX8446);
  dff DFF_1207(CK,WX8449,WX8448);
  dff DFF_1208(CK,WX8451,WX8450);
  dff DFF_1209(CK,WX8453,WX8452);
  dff DFF_1210(CK,WX8455,WX8454);
  dff DFF_1211(CK,WX8457,WX8456);
  dff DFF_1212(CK,WX8459,WX8458);
  dff DFF_1213(CK,WX8461,WX8460);
  dff DFF_1214(CK,WX8463,WX8462);
  dff DFF_1215(CK,WX8465,WX8464);
  dff DFF_1216(CK,WX8467,WX8466);
  dff DFF_1217(CK,WX8469,WX8468);
  dff DFF_1218(CK,WX8471,WX8470);
  dff DFF_1219(CK,WX8473,WX8472);
  dff DFF_1220(CK,WX8475,WX8474);
  dff DFF_1221(CK,WX8477,WX8476);
  dff DFF_1222(CK,WX8479,WX8478);
  dff DFF_1223(CK,WX8481,WX8480);
  dff DFF_1224(CK,WX8483,WX8482);
  dff DFF_1225(CK,WX8485,WX8484);
  dff DFF_1226(CK,WX8487,WX8486);
  dff DFF_1227(CK,WX8489,WX8488);
  dff DFF_1228(CK,WX8491,WX8490);
  dff DFF_1229(CK,WX8493,WX8492);
  dff DFF_1230(CK,WX8495,WX8494);
  dff DFF_1231(CK,WX8497,WX8496);
  dff DFF_1232(CK,WX8499,WX8498);
  dff DFF_1233(CK,WX8501,WX8500);
  dff DFF_1234(CK,WX8503,WX8502);
  dff DFF_1235(CK,WX8505,WX8504);
  dff DFF_1236(CK,WX8507,WX8506);
  dff DFF_1237(CK,WX8509,WX8508);
  dff DFF_1238(CK,WX8511,WX8510);
  dff DFF_1239(CK,WX8513,WX8512);
  dff DFF_1240(CK,WX8515,WX8514);
  dff DFF_1241(CK,WX8517,WX8516);
  dff DFF_1242(CK,WX8519,WX8518);
  dff DFF_1243(CK,WX8521,WX8520);
  dff DFF_1244(CK,WX8523,WX8522);
  dff DFF_1245(CK,WX8525,WX8524);
  dff DFF_1246(CK,WX8527,WX8526);
  dff DFF_1247(CK,WX8529,WX8528);
  dff DFF_1248(CK,WX8531,WX8530);
  dff DFF_1249(CK,WX8533,WX8532);
  dff DFF_1250(CK,WX8535,WX8534);
  dff DFF_1251(CK,WX8537,WX8536);
  dff DFF_1252(CK,WX8539,WX8538);
  dff DFF_1253(CK,WX8541,WX8540);
  dff DFF_1254(CK,WX8543,WX8542);
  dff DFF_1255(CK,WX8545,WX8544);
  dff DFF_1256(CK,WX8547,WX8546);
  dff DFF_1257(CK,WX8549,WX8548);
  dff DFF_1258(CK,WX8551,WX8550);
  dff DFF_1259(CK,WX8553,WX8552);
  dff DFF_1260(CK,WX8555,WX8554);
  dff DFF_1261(CK,WX8557,WX8556);
  dff DFF_1262(CK,WX8559,WX8558);
  dff DFF_1263(CK,WX8561,WX8560);
  dff DFF_1264(CK,WX8563,WX8562);
  dff DFF_1265(CK,WX8565,WX8564);
  dff DFF_1266(CK,WX8567,WX8566);
  dff DFF_1267(CK,WX8569,WX8568);
  dff DFF_1268(CK,WX8571,WX8570);
  dff DFF_1269(CK,WX8573,WX8572);
  dff DFF_1270(CK,WX8575,WX8574);
  dff DFF_1271(CK,WX8577,WX8576);
  dff DFF_1272(CK,WX8579,WX8578);
  dff DFF_1273(CK,WX8581,WX8580);
  dff DFF_1274(CK,WX8583,WX8582);
  dff DFF_1275(CK,WX8585,WX8584);
  dff DFF_1276(CK,WX8587,WX8586);
  dff DFF_1277(CK,WX8589,WX8588);
  dff DFF_1278(CK,WX8591,WX8590);
  dff DFF_1279(CK,WX8593,WX8592);
  dff DFF_1280(CK,WX8595,WX8594);
  dff DFF_1281(CK,WX8597,WX8596);
  dff DFF_1282(CK,WX8599,WX8598);
  dff DFF_1283(CK,WX8601,WX8600);
  dff DFF_1284(CK,WX8603,WX8602);
  dff DFF_1285(CK,WX8605,WX8604);
  dff DFF_1286(CK,WX8607,WX8606);
  dff DFF_1287(CK,WX8609,WX8608);
  dff DFF_1288(CK,WX8611,WX8610);
  dff DFF_1289(CK,WX8613,WX8612);
  dff DFF_1290(CK,WX8615,WX8614);
  dff DFF_1291(CK,WX8617,WX8616);
  dff DFF_1292(CK,WX8619,WX8618);
  dff DFF_1293(CK,WX8621,WX8620);
  dff DFF_1294(CK,WX8623,WX8622);
  dff DFF_1295(CK,WX8625,WX8624);
  dff DFF_1296(CK,WX8627,WX8626);
  dff DFF_1297(CK,WX8629,WX8628);
  dff DFF_1298(CK,WX8631,WX8630);
  dff DFF_1299(CK,WX8633,WX8632);
  dff DFF_1300(CK,WX8635,WX8634);
  dff DFF_1301(CK,WX8637,WX8636);
  dff DFF_1302(CK,WX8639,WX8638);
  dff DFF_1303(CK,WX8641,WX8640);
  dff DFF_1304(CK,WX8643,WX8642);
  dff DFF_1305(CK,WX8645,WX8644);
  dff DFF_1306(CK,WX8647,WX8646);
  dff DFF_1307(CK,WX8649,WX8648);
  dff DFF_1308(CK,WX8651,WX8650);
  dff DFF_1309(CK,WX8653,WX8652);
  dff DFF_1310(CK,WX8655,WX8654);
  dff DFF_1311(CK,WX8657,WX8656);
  dff DFF_1312(CK,CRC_OUT_3_0,WX9022);
  dff DFF_1313(CK,CRC_OUT_3_1,WX9024);
  dff DFF_1314(CK,CRC_OUT_3_2,WX9026);
  dff DFF_1315(CK,CRC_OUT_3_3,WX9028);
  dff DFF_1316(CK,CRC_OUT_3_4,WX9030);
  dff DFF_1317(CK,CRC_OUT_3_5,WX9032);
  dff DFF_1318(CK,CRC_OUT_3_6,WX9034);
  dff DFF_1319(CK,CRC_OUT_3_7,WX9036);
  dff DFF_1320(CK,CRC_OUT_3_8,WX9038);
  dff DFF_1321(CK,CRC_OUT_3_9,WX9040);
  dff DFF_1322(CK,CRC_OUT_3_10,WX9042);
  dff DFF_1323(CK,CRC_OUT_3_11,WX9044);
  dff DFF_1324(CK,CRC_OUT_3_12,WX9046);
  dff DFF_1325(CK,CRC_OUT_3_13,WX9048);
  dff DFF_1326(CK,CRC_OUT_3_14,WX9050);
  dff DFF_1327(CK,CRC_OUT_3_15,WX9052);
  dff DFF_1328(CK,CRC_OUT_3_16,WX9054);
  dff DFF_1329(CK,CRC_OUT_3_17,WX9056);
  dff DFF_1330(CK,CRC_OUT_3_18,WX9058);
  dff DFF_1331(CK,CRC_OUT_3_19,WX9060);
  dff DFF_1332(CK,CRC_OUT_3_20,WX9062);
  dff DFF_1333(CK,CRC_OUT_3_21,WX9064);
  dff DFF_1334(CK,CRC_OUT_3_22,WX9066);
  dff DFF_1335(CK,CRC_OUT_3_23,WX9068);
  dff DFF_1336(CK,CRC_OUT_3_24,WX9070);
  dff DFF_1337(CK,CRC_OUT_3_25,WX9072);
  dff DFF_1338(CK,CRC_OUT_3_26,WX9074);
  dff DFF_1339(CK,CRC_OUT_3_27,WX9076);
  dff DFF_1340(CK,CRC_OUT_3_28,WX9078);
  dff DFF_1341(CK,CRC_OUT_3_29,WX9080);
  dff DFF_1342(CK,CRC_OUT_3_30,WX9082);
  dff DFF_1343(CK,CRC_OUT_3_31,WX9084);
  dff DFF_1344(CK,WX9536,WX9535);
  dff DFF_1345(CK,WX9538,WX9537);
  dff DFF_1346(CK,WX9540,WX9539);
  dff DFF_1347(CK,WX9542,WX9541);
  dff DFF_1348(CK,WX9544,WX9543);
  dff DFF_1349(CK,WX9546,WX9545);
  dff DFF_1350(CK,WX9548,WX9547);
  dff DFF_1351(CK,WX9550,WX9549);
  dff DFF_1352(CK,WX9552,WX9551);
  dff DFF_1353(CK,WX9554,WX9553);
  dff DFF_1354(CK,WX9556,WX9555);
  dff DFF_1355(CK,WX9558,WX9557);
  dff DFF_1356(CK,WX9560,WX9559);
  dff DFF_1357(CK,WX9562,WX9561);
  dff DFF_1358(CK,WX9564,WX9563);
  dff DFF_1359(CK,WX9566,WX9565);
  dff DFF_1360(CK,WX9568,WX9567);
  dff DFF_1361(CK,WX9570,WX9569);
  dff DFF_1362(CK,WX9572,WX9571);
  dff DFF_1363(CK,WX9574,WX9573);
  dff DFF_1364(CK,WX9576,WX9575);
  dff DFF_1365(CK,WX9578,WX9577);
  dff DFF_1366(CK,WX9580,WX9579);
  dff DFF_1367(CK,WX9582,WX9581);
  dff DFF_1368(CK,WX9584,WX9583);
  dff DFF_1369(CK,WX9586,WX9585);
  dff DFF_1370(CK,WX9588,WX9587);
  dff DFF_1371(CK,WX9590,WX9589);
  dff DFF_1372(CK,WX9592,WX9591);
  dff DFF_1373(CK,WX9594,WX9593);
  dff DFF_1374(CK,WX9596,WX9595);
  dff DFF_1375(CK,WX9598,WX9597);
  dff DFF_1376(CK,WX9696,WX9695);
  dff DFF_1377(CK,WX9698,WX9697);
  dff DFF_1378(CK,WX9700,WX9699);
  dff DFF_1379(CK,WX9702,WX9701);
  dff DFF_1380(CK,WX9704,WX9703);
  dff DFF_1381(CK,WX9706,WX9705);
  dff DFF_1382(CK,WX9708,WX9707);
  dff DFF_1383(CK,WX9710,WX9709);
  dff DFF_1384(CK,WX9712,WX9711);
  dff DFF_1385(CK,WX9714,WX9713);
  dff DFF_1386(CK,WX9716,WX9715);
  dff DFF_1387(CK,WX9718,WX9717);
  dff DFF_1388(CK,WX9720,WX9719);
  dff DFF_1389(CK,WX9722,WX9721);
  dff DFF_1390(CK,WX9724,WX9723);
  dff DFF_1391(CK,WX9726,WX9725);
  dff DFF_1392(CK,WX9728,WX9727);
  dff DFF_1393(CK,WX9730,WX9729);
  dff DFF_1394(CK,WX9732,WX9731);
  dff DFF_1395(CK,WX9734,WX9733);
  dff DFF_1396(CK,WX9736,WX9735);
  dff DFF_1397(CK,WX9738,WX9737);
  dff DFF_1398(CK,WX9740,WX9739);
  dff DFF_1399(CK,WX9742,WX9741);
  dff DFF_1400(CK,WX9744,WX9743);
  dff DFF_1401(CK,WX9746,WX9745);
  dff DFF_1402(CK,WX9748,WX9747);
  dff DFF_1403(CK,WX9750,WX9749);
  dff DFF_1404(CK,WX9752,WX9751);
  dff DFF_1405(CK,WX9754,WX9753);
  dff DFF_1406(CK,WX9756,WX9755);
  dff DFF_1407(CK,WX9758,WX9757);
  dff DFF_1408(CK,WX9760,WX9759);
  dff DFF_1409(CK,WX9762,WX9761);
  dff DFF_1410(CK,WX9764,WX9763);
  dff DFF_1411(CK,WX9766,WX9765);
  dff DFF_1412(CK,WX9768,WX9767);
  dff DFF_1413(CK,WX9770,WX9769);
  dff DFF_1414(CK,WX9772,WX9771);
  dff DFF_1415(CK,WX9774,WX9773);
  dff DFF_1416(CK,WX9776,WX9775);
  dff DFF_1417(CK,WX9778,WX9777);
  dff DFF_1418(CK,WX9780,WX9779);
  dff DFF_1419(CK,WX9782,WX9781);
  dff DFF_1420(CK,WX9784,WX9783);
  dff DFF_1421(CK,WX9786,WX9785);
  dff DFF_1422(CK,WX9788,WX9787);
  dff DFF_1423(CK,WX9790,WX9789);
  dff DFF_1424(CK,WX9792,WX9791);
  dff DFF_1425(CK,WX9794,WX9793);
  dff DFF_1426(CK,WX9796,WX9795);
  dff DFF_1427(CK,WX9798,WX9797);
  dff DFF_1428(CK,WX9800,WX9799);
  dff DFF_1429(CK,WX9802,WX9801);
  dff DFF_1430(CK,WX9804,WX9803);
  dff DFF_1431(CK,WX9806,WX9805);
  dff DFF_1432(CK,WX9808,WX9807);
  dff DFF_1433(CK,WX9810,WX9809);
  dff DFF_1434(CK,WX9812,WX9811);
  dff DFF_1435(CK,WX9814,WX9813);
  dff DFF_1436(CK,WX9816,WX9815);
  dff DFF_1437(CK,WX9818,WX9817);
  dff DFF_1438(CK,WX9820,WX9819);
  dff DFF_1439(CK,WX9822,WX9821);
  dff DFF_1440(CK,WX9824,WX9823);
  dff DFF_1441(CK,WX9826,WX9825);
  dff DFF_1442(CK,WX9828,WX9827);
  dff DFF_1443(CK,WX9830,WX9829);
  dff DFF_1444(CK,WX9832,WX9831);
  dff DFF_1445(CK,WX9834,WX9833);
  dff DFF_1446(CK,WX9836,WX9835);
  dff DFF_1447(CK,WX9838,WX9837);
  dff DFF_1448(CK,WX9840,WX9839);
  dff DFF_1449(CK,WX9842,WX9841);
  dff DFF_1450(CK,WX9844,WX9843);
  dff DFF_1451(CK,WX9846,WX9845);
  dff DFF_1452(CK,WX9848,WX9847);
  dff DFF_1453(CK,WX9850,WX9849);
  dff DFF_1454(CK,WX9852,WX9851);
  dff DFF_1455(CK,WX9854,WX9853);
  dff DFF_1456(CK,WX9856,WX9855);
  dff DFF_1457(CK,WX9858,WX9857);
  dff DFF_1458(CK,WX9860,WX9859);
  dff DFF_1459(CK,WX9862,WX9861);
  dff DFF_1460(CK,WX9864,WX9863);
  dff DFF_1461(CK,WX9866,WX9865);
  dff DFF_1462(CK,WX9868,WX9867);
  dff DFF_1463(CK,WX9870,WX9869);
  dff DFF_1464(CK,WX9872,WX9871);
  dff DFF_1465(CK,WX9874,WX9873);
  dff DFF_1466(CK,WX9876,WX9875);
  dff DFF_1467(CK,WX9878,WX9877);
  dff DFF_1468(CK,WX9880,WX9879);
  dff DFF_1469(CK,WX9882,WX9881);
  dff DFF_1470(CK,WX9884,WX9883);
  dff DFF_1471(CK,WX9886,WX9885);
  dff DFF_1472(CK,WX9888,WX9887);
  dff DFF_1473(CK,WX9890,WX9889);
  dff DFF_1474(CK,WX9892,WX9891);
  dff DFF_1475(CK,WX9894,WX9893);
  dff DFF_1476(CK,WX9896,WX9895);
  dff DFF_1477(CK,WX9898,WX9897);
  dff DFF_1478(CK,WX9900,WX9899);
  dff DFF_1479(CK,WX9902,WX9901);
  dff DFF_1480(CK,WX9904,WX9903);
  dff DFF_1481(CK,WX9906,WX9905);
  dff DFF_1482(CK,WX9908,WX9907);
  dff DFF_1483(CK,WX9910,WX9909);
  dff DFF_1484(CK,WX9912,WX9911);
  dff DFF_1485(CK,WX9914,WX9913);
  dff DFF_1486(CK,WX9916,WX9915);
  dff DFF_1487(CK,WX9918,WX9917);
  dff DFF_1488(CK,WX9920,WX9919);
  dff DFF_1489(CK,WX9922,WX9921);
  dff DFF_1490(CK,WX9924,WX9923);
  dff DFF_1491(CK,WX9926,WX9925);
  dff DFF_1492(CK,WX9928,WX9927);
  dff DFF_1493(CK,WX9930,WX9929);
  dff DFF_1494(CK,WX9932,WX9931);
  dff DFF_1495(CK,WX9934,WX9933);
  dff DFF_1496(CK,WX9936,WX9935);
  dff DFF_1497(CK,WX9938,WX9937);
  dff DFF_1498(CK,WX9940,WX9939);
  dff DFF_1499(CK,WX9942,WX9941);
  dff DFF_1500(CK,WX9944,WX9943);
  dff DFF_1501(CK,WX9946,WX9945);
  dff DFF_1502(CK,WX9948,WX9947);
  dff DFF_1503(CK,WX9950,WX9949);
  dff DFF_1504(CK,CRC_OUT_2_0,WX10315);
  dff DFF_1505(CK,CRC_OUT_2_1,WX10317);
  dff DFF_1506(CK,CRC_OUT_2_2,WX10319);
  dff DFF_1507(CK,CRC_OUT_2_3,WX10321);
  dff DFF_1508(CK,CRC_OUT_2_4,WX10323);
  dff DFF_1509(CK,CRC_OUT_2_5,WX10325);
  dff DFF_1510(CK,CRC_OUT_2_6,WX10327);
  dff DFF_1511(CK,CRC_OUT_2_7,WX10329);
  dff DFF_1512(CK,CRC_OUT_2_8,WX10331);
  dff DFF_1513(CK,CRC_OUT_2_9,WX10333);
  dff DFF_1514(CK,CRC_OUT_2_10,WX10335);
  dff DFF_1515(CK,CRC_OUT_2_11,WX10337);
  dff DFF_1516(CK,CRC_OUT_2_12,WX10339);
  dff DFF_1517(CK,CRC_OUT_2_13,WX10341);
  dff DFF_1518(CK,CRC_OUT_2_14,WX10343);
  dff DFF_1519(CK,CRC_OUT_2_15,WX10345);
  dff DFF_1520(CK,CRC_OUT_2_16,WX10347);
  dff DFF_1521(CK,CRC_OUT_2_17,WX10349);
  dff DFF_1522(CK,CRC_OUT_2_18,WX10351);
  dff DFF_1523(CK,CRC_OUT_2_19,WX10353);
  dff DFF_1524(CK,CRC_OUT_2_20,WX10355);
  dff DFF_1525(CK,CRC_OUT_2_21,WX10357);
  dff DFF_1526(CK,CRC_OUT_2_22,WX10359);
  dff DFF_1527(CK,CRC_OUT_2_23,WX10361);
  dff DFF_1528(CK,CRC_OUT_2_24,WX10363);
  dff DFF_1529(CK,CRC_OUT_2_25,WX10365);
  dff DFF_1530(CK,CRC_OUT_2_26,WX10367);
  dff DFF_1531(CK,CRC_OUT_2_27,WX10369);
  dff DFF_1532(CK,CRC_OUT_2_28,WX10371);
  dff DFF_1533(CK,CRC_OUT_2_29,WX10373);
  dff DFF_1534(CK,CRC_OUT_2_30,WX10375);
  dff DFF_1535(CK,CRC_OUT_2_31,WX10377);
  dff DFF_1536(CK,WX10829,WX10828);
  dff DFF_1537(CK,WX10831,WX10830);
  dff DFF_1538(CK,WX10833,WX10832);
  dff DFF_1539(CK,WX10835,WX10834);
  dff DFF_1540(CK,WX10837,WX10836);
  dff DFF_1541(CK,WX10839,WX10838);
  dff DFF_1542(CK,WX10841,WX10840);
  dff DFF_1543(CK,WX10843,WX10842);
  dff DFF_1544(CK,WX10845,WX10844);
  dff DFF_1545(CK,WX10847,WX10846);
  dff DFF_1546(CK,WX10849,WX10848);
  dff DFF_1547(CK,WX10851,WX10850);
  dff DFF_1548(CK,WX10853,WX10852);
  dff DFF_1549(CK,WX10855,WX10854);
  dff DFF_1550(CK,WX10857,WX10856);
  dff DFF_1551(CK,WX10859,WX10858);
  dff DFF_1552(CK,WX10861,WX10860);
  dff DFF_1553(CK,WX10863,WX10862);
  dff DFF_1554(CK,WX10865,WX10864);
  dff DFF_1555(CK,WX10867,WX10866);
  dff DFF_1556(CK,WX10869,WX10868);
  dff DFF_1557(CK,WX10871,WX10870);
  dff DFF_1558(CK,WX10873,WX10872);
  dff DFF_1559(CK,WX10875,WX10874);
  dff DFF_1560(CK,WX10877,WX10876);
  dff DFF_1561(CK,WX10879,WX10878);
  dff DFF_1562(CK,WX10881,WX10880);
  dff DFF_1563(CK,WX10883,WX10882);
  dff DFF_1564(CK,WX10885,WX10884);
  dff DFF_1565(CK,WX10887,WX10886);
  dff DFF_1566(CK,WX10889,WX10888);
  dff DFF_1567(CK,WX10891,WX10890);
  dff DFF_1568(CK,WX10989,WX10988);
  dff DFF_1569(CK,WX10991,WX10990);
  dff DFF_1570(CK,WX10993,WX10992);
  dff DFF_1571(CK,WX10995,WX10994);
  dff DFF_1572(CK,WX10997,WX10996);
  dff DFF_1573(CK,WX10999,WX10998);
  dff DFF_1574(CK,WX11001,WX11000);
  dff DFF_1575(CK,WX11003,WX11002);
  dff DFF_1576(CK,WX11005,WX11004);
  dff DFF_1577(CK,WX11007,WX11006);
  dff DFF_1578(CK,WX11009,WX11008);
  dff DFF_1579(CK,WX11011,WX11010);
  dff DFF_1580(CK,WX11013,WX11012);
  dff DFF_1581(CK,WX11015,WX11014);
  dff DFF_1582(CK,WX11017,WX11016);
  dff DFF_1583(CK,WX11019,WX11018);
  dff DFF_1584(CK,WX11021,WX11020);
  dff DFF_1585(CK,WX11023,WX11022);
  dff DFF_1586(CK,WX11025,WX11024);
  dff DFF_1587(CK,WX11027,WX11026);
  dff DFF_1588(CK,WX11029,WX11028);
  dff DFF_1589(CK,WX11031,WX11030);
  dff DFF_1590(CK,WX11033,WX11032);
  dff DFF_1591(CK,WX11035,WX11034);
  dff DFF_1592(CK,WX11037,WX11036);
  dff DFF_1593(CK,WX11039,WX11038);
  dff DFF_1594(CK,WX11041,WX11040);
  dff DFF_1595(CK,WX11043,WX11042);
  dff DFF_1596(CK,WX11045,WX11044);
  dff DFF_1597(CK,WX11047,WX11046);
  dff DFF_1598(CK,WX11049,WX11048);
  dff DFF_1599(CK,WX11051,WX11050);
  dff DFF_1600(CK,WX11053,WX11052);
  dff DFF_1601(CK,WX11055,WX11054);
  dff DFF_1602(CK,WX11057,WX11056);
  dff DFF_1603(CK,WX11059,WX11058);
  dff DFF_1604(CK,WX11061,WX11060);
  dff DFF_1605(CK,WX11063,WX11062);
  dff DFF_1606(CK,WX11065,WX11064);
  dff DFF_1607(CK,WX11067,WX11066);
  dff DFF_1608(CK,WX11069,WX11068);
  dff DFF_1609(CK,WX11071,WX11070);
  dff DFF_1610(CK,WX11073,WX11072);
  dff DFF_1611(CK,WX11075,WX11074);
  dff DFF_1612(CK,WX11077,WX11076);
  dff DFF_1613(CK,WX11079,WX11078);
  dff DFF_1614(CK,WX11081,WX11080);
  dff DFF_1615(CK,WX11083,WX11082);
  dff DFF_1616(CK,WX11085,WX11084);
  dff DFF_1617(CK,WX11087,WX11086);
  dff DFF_1618(CK,WX11089,WX11088);
  dff DFF_1619(CK,WX11091,WX11090);
  dff DFF_1620(CK,WX11093,WX11092);
  dff DFF_1621(CK,WX11095,WX11094);
  dff DFF_1622(CK,WX11097,WX11096);
  dff DFF_1623(CK,WX11099,WX11098);
  dff DFF_1624(CK,WX11101,WX11100);
  dff DFF_1625(CK,WX11103,WX11102);
  dff DFF_1626(CK,WX11105,WX11104);
  dff DFF_1627(CK,WX11107,WX11106);
  dff DFF_1628(CK,WX11109,WX11108);
  dff DFF_1629(CK,WX11111,WX11110);
  dff DFF_1630(CK,WX11113,WX11112);
  dff DFF_1631(CK,WX11115,WX11114);
  dff DFF_1632(CK,WX11117,WX11116);
  dff DFF_1633(CK,WX11119,WX11118);
  dff DFF_1634(CK,WX11121,WX11120);
  dff DFF_1635(CK,WX11123,WX11122);
  dff DFF_1636(CK,WX11125,WX11124);
  dff DFF_1637(CK,WX11127,WX11126);
  dff DFF_1638(CK,WX11129,WX11128);
  dff DFF_1639(CK,WX11131,WX11130);
  dff DFF_1640(CK,WX11133,WX11132);
  dff DFF_1641(CK,WX11135,WX11134);
  dff DFF_1642(CK,WX11137,WX11136);
  dff DFF_1643(CK,WX11139,WX11138);
  dff DFF_1644(CK,WX11141,WX11140);
  dff DFF_1645(CK,WX11143,WX11142);
  dff DFF_1646(CK,WX11145,WX11144);
  dff DFF_1647(CK,WX11147,WX11146);
  dff DFF_1648(CK,WX11149,WX11148);
  dff DFF_1649(CK,WX11151,WX11150);
  dff DFF_1650(CK,WX11153,WX11152);
  dff DFF_1651(CK,WX11155,WX11154);
  dff DFF_1652(CK,WX11157,WX11156);
  dff DFF_1653(CK,WX11159,WX11158);
  dff DFF_1654(CK,WX11161,WX11160);
  dff DFF_1655(CK,WX11163,WX11162);
  dff DFF_1656(CK,WX11165,WX11164);
  dff DFF_1657(CK,WX11167,WX11166);
  dff DFF_1658(CK,WX11169,WX11168);
  dff DFF_1659(CK,WX11171,WX11170);
  dff DFF_1660(CK,WX11173,WX11172);
  dff DFF_1661(CK,WX11175,WX11174);
  dff DFF_1662(CK,WX11177,WX11176);
  dff DFF_1663(CK,WX11179,WX11178);
  dff DFF_1664(CK,WX11181,WX11180);
  dff DFF_1665(CK,WX11183,WX11182);
  dff DFF_1666(CK,WX11185,WX11184);
  dff DFF_1667(CK,WX11187,WX11186);
  dff DFF_1668(CK,WX11189,WX11188);
  dff DFF_1669(CK,WX11191,WX11190);
  dff DFF_1670(CK,WX11193,WX11192);
  dff DFF_1671(CK,WX11195,WX11194);
  dff DFF_1672(CK,WX11197,WX11196);
  dff DFF_1673(CK,WX11199,WX11198);
  dff DFF_1674(CK,WX11201,WX11200);
  dff DFF_1675(CK,WX11203,WX11202);
  dff DFF_1676(CK,WX11205,WX11204);
  dff DFF_1677(CK,WX11207,WX11206);
  dff DFF_1678(CK,WX11209,WX11208);
  dff DFF_1679(CK,WX11211,WX11210);
  dff DFF_1680(CK,WX11213,WX11212);
  dff DFF_1681(CK,WX11215,WX11214);
  dff DFF_1682(CK,WX11217,WX11216);
  dff DFF_1683(CK,WX11219,WX11218);
  dff DFF_1684(CK,WX11221,WX11220);
  dff DFF_1685(CK,WX11223,WX11222);
  dff DFF_1686(CK,WX11225,WX11224);
  dff DFF_1687(CK,WX11227,WX11226);
  dff DFF_1688(CK,WX11229,WX11228);
  dff DFF_1689(CK,WX11231,WX11230);
  dff DFF_1690(CK,WX11233,WX11232);
  dff DFF_1691(CK,WX11235,WX11234);
  dff DFF_1692(CK,WX11237,WX11236);
  dff DFF_1693(CK,WX11239,WX11238);
  dff DFF_1694(CK,WX11241,WX11240);
  dff DFF_1695(CK,WX11243,WX11242);
  dff DFF_1696(CK,CRC_OUT_1_0,WX11608);
  dff DFF_1697(CK,CRC_OUT_1_1,WX11610);
  dff DFF_1698(CK,CRC_OUT_1_2,WX11612);
  dff DFF_1699(CK,CRC_OUT_1_3,WX11614);
  dff DFF_1700(CK,CRC_OUT_1_4,WX11616);
  dff DFF_1701(CK,CRC_OUT_1_5,WX11618);
  dff DFF_1702(CK,CRC_OUT_1_6,WX11620);
  dff DFF_1703(CK,CRC_OUT_1_7,WX11622);
  dff DFF_1704(CK,CRC_OUT_1_8,WX11624);
  dff DFF_1705(CK,CRC_OUT_1_9,WX11626);
  dff DFF_1706(CK,CRC_OUT_1_10,WX11628);
  dff DFF_1707(CK,CRC_OUT_1_11,WX11630);
  dff DFF_1708(CK,CRC_OUT_1_12,WX11632);
  dff DFF_1709(CK,CRC_OUT_1_13,WX11634);
  dff DFF_1710(CK,CRC_OUT_1_14,WX11636);
  dff DFF_1711(CK,CRC_OUT_1_15,WX11638);
  dff DFF_1712(CK,CRC_OUT_1_16,WX11640);
  dff DFF_1713(CK,CRC_OUT_1_17,WX11642);
  dff DFF_1714(CK,CRC_OUT_1_18,WX11644);
  dff DFF_1715(CK,CRC_OUT_1_19,WX11646);
  dff DFF_1716(CK,CRC_OUT_1_20,WX11648);
  dff DFF_1717(CK,CRC_OUT_1_21,WX11650);
  dff DFF_1718(CK,CRC_OUT_1_22,WX11652);
  dff DFF_1719(CK,CRC_OUT_1_23,WX11654);
  dff DFF_1720(CK,CRC_OUT_1_24,WX11656);
  dff DFF_1721(CK,CRC_OUT_1_25,WX11658);
  dff DFF_1722(CK,CRC_OUT_1_26,WX11660);
  dff DFF_1723(CK,CRC_OUT_1_27,WX11662);
  dff DFF_1724(CK,CRC_OUT_1_28,WX11664);
  dff DFF_1725(CK,CRC_OUT_1_29,WX11666);
  dff DFF_1726(CK,CRC_OUT_1_30,WX11668);
  dff DFF_1727(CK,CRC_OUT_1_31,WX11670);
  not NOT_0(WX37,WX1003);
  not NOT_1(WX41,WX1004);
  not NOT_2(WX45,WX1004);
  not NOT_3(WX47,WX38);
  not NOT_4(WX48,WX47);
  not NOT_5(WX51,WX1003);
  not NOT_6(WX55,WX1004);
  not NOT_7(WX59,WX1004);
  not NOT_8(WX61,WX52);
  not NOT_9(WX62,WX61);
  not NOT_10(WX65,WX1003);
  not NOT_11(WX69,WX1004);
  not NOT_12(WX73,WX1004);
  not NOT_13(WX75,WX66);
  not NOT_14(WX76,WX75);
  not NOT_15(WX79,WX1003);
  not NOT_16(WX83,WX1004);
  not NOT_17(WX87,WX1004);
  not NOT_18(WX89,WX80);
  not NOT_19(WX90,WX89);
  not NOT_20(WX93,WX1003);
  not NOT_21(WX97,WX1004);
  not NOT_22(WX101,WX1004);
  not NOT_23(WX103,WX94);
  not NOT_24(WX104,WX103);
  not NOT_25(WX107,WX1003);
  not NOT_26(WX111,WX1004);
  not NOT_27(WX115,WX1004);
  not NOT_28(WX117,WX108);
  not NOT_29(WX118,WX117);
  not NOT_30(WX121,WX1003);
  not NOT_31(WX125,WX1004);
  not NOT_32(WX129,WX1004);
  not NOT_33(WX131,WX122);
  not NOT_34(WX132,WX131);
  not NOT_35(WX135,WX1003);
  not NOT_36(WX139,WX1004);
  not NOT_37(WX143,WX1004);
  not NOT_38(WX145,WX136);
  not NOT_39(WX146,WX145);
  not NOT_40(WX149,WX1003);
  not NOT_41(WX153,WX1004);
  not NOT_42(WX157,WX1004);
  not NOT_43(WX159,WX150);
  not NOT_44(WX160,WX159);
  not NOT_45(WX163,WX1003);
  not NOT_46(WX167,WX1004);
  not NOT_47(WX171,WX1004);
  not NOT_48(WX173,WX164);
  not NOT_49(WX174,WX173);
  not NOT_50(WX177,WX1003);
  not NOT_51(WX181,WX1004);
  not NOT_52(WX185,WX1004);
  not NOT_53(WX187,WX178);
  not NOT_54(WX188,WX187);
  not NOT_55(WX191,WX1003);
  not NOT_56(WX195,WX1004);
  not NOT_57(WX199,WX1004);
  not NOT_58(WX201,WX192);
  not NOT_59(WX202,WX201);
  not NOT_60(WX205,WX1003);
  not NOT_61(WX209,WX1004);
  not NOT_62(WX213,WX1004);
  not NOT_63(WX215,WX206);
  not NOT_64(WX216,WX215);
  not NOT_65(WX219,WX1003);
  not NOT_66(WX223,WX1004);
  not NOT_67(WX227,WX1004);
  not NOT_68(WX229,WX220);
  not NOT_69(WX230,WX229);
  not NOT_70(WX233,WX1003);
  not NOT_71(WX237,WX1004);
  not NOT_72(WX241,WX1004);
  not NOT_73(WX243,WX234);
  not NOT_74(WX244,WX243);
  not NOT_75(WX247,WX1003);
  not NOT_76(WX251,WX1004);
  not NOT_77(WX255,WX1004);
  not NOT_78(WX257,WX248);
  not NOT_79(WX258,WX257);
  not NOT_80(WX261,WX1003);
  not NOT_81(WX265,WX1004);
  not NOT_82(WX269,WX1004);
  not NOT_83(WX271,WX262);
  not NOT_84(WX272,WX271);
  not NOT_85(WX275,WX1003);
  not NOT_86(WX279,WX1004);
  not NOT_87(WX283,WX1004);
  not NOT_88(WX285,WX276);
  not NOT_89(WX286,WX285);
  not NOT_90(WX289,WX1003);
  not NOT_91(WX293,WX1004);
  not NOT_92(WX297,WX1004);
  not NOT_93(WX299,WX290);
  not NOT_94(WX300,WX299);
  not NOT_95(WX303,WX1003);
  not NOT_96(WX307,WX1004);
  not NOT_97(WX311,WX1004);
  not NOT_98(WX313,WX304);
  not NOT_99(WX314,WX313);
  not NOT_100(WX317,WX1003);
  not NOT_101(WX321,WX1004);
  not NOT_102(WX325,WX1004);
  not NOT_103(WX327,WX318);
  not NOT_104(WX328,WX327);
  not NOT_105(WX331,WX1003);
  not NOT_106(WX335,WX1004);
  not NOT_107(WX339,WX1004);
  not NOT_108(WX341,WX332);
  not NOT_109(WX342,WX341);
  not NOT_110(WX345,WX1003);
  not NOT_111(WX349,WX1004);
  not NOT_112(WX353,WX1004);
  not NOT_113(WX355,WX346);
  not NOT_114(WX356,WX355);
  not NOT_115(WX359,WX1003);
  not NOT_116(WX363,WX1004);
  not NOT_117(WX367,WX1004);
  not NOT_118(WX369,WX360);
  not NOT_119(WX370,WX369);
  not NOT_120(WX373,WX1003);
  not NOT_121(WX377,WX1004);
  not NOT_122(WX381,WX1004);
  not NOT_123(WX383,WX374);
  not NOT_124(WX384,WX383);
  not NOT_125(WX387,WX1003);
  not NOT_126(WX391,WX1004);
  not NOT_127(WX395,WX1004);
  not NOT_128(WX397,WX388);
  not NOT_129(WX398,WX397);
  not NOT_130(WX401,WX1003);
  not NOT_131(WX405,WX1004);
  not NOT_132(WX409,WX1004);
  not NOT_133(WX411,WX402);
  not NOT_134(WX412,WX411);
  not NOT_135(WX415,WX1003);
  not NOT_136(WX419,WX1004);
  not NOT_137(WX423,WX1004);
  not NOT_138(WX425,WX416);
  not NOT_139(WX426,WX425);
  not NOT_140(WX429,WX1003);
  not NOT_141(WX433,WX1004);
  not NOT_142(WX437,WX1004);
  not NOT_143(WX439,WX430);
  not NOT_144(WX440,WX439);
  not NOT_145(WX443,WX1003);
  not NOT_146(WX447,WX1004);
  not NOT_147(WX451,WX1004);
  not NOT_148(WX453,WX444);
  not NOT_149(WX454,WX453);
  not NOT_150(WX457,WX1003);
  not NOT_151(WX461,WX1004);
  not NOT_152(WX465,WX1004);
  not NOT_153(WX467,WX458);
  not NOT_154(WX468,WX467);
  not NOT_155(WX471,WX1003);
  not NOT_156(WX475,WX1004);
  not NOT_157(WX479,WX1004);
  not NOT_158(WX481,WX472);
  not NOT_159(WX482,WX481);
  not NOT_160(WX483,WX485);
  not NOT_161(WX548,WX965);
  not NOT_162(WX549,WX967);
  not NOT_163(WX550,WX969);
  not NOT_164(WX551,WX971);
  not NOT_165(WX552,WX973);
  not NOT_166(WX553,WX975);
  not NOT_167(WX554,WX977);
  not NOT_168(WX555,WX979);
  not NOT_169(WX556,WX981);
  not NOT_170(WX557,WX983);
  not NOT_171(WX558,WX985);
  not NOT_172(WX559,WX987);
  not NOT_173(WX560,WX989);
  not NOT_174(WX561,WX991);
  not NOT_175(WX562,WX993);
  not NOT_176(WX563,WX995);
  not NOT_177(WX564,WX933);
  not NOT_178(WX565,WX935);
  not NOT_179(WX566,WX937);
  not NOT_180(WX567,WX939);
  not NOT_181(WX568,WX941);
  not NOT_182(WX569,WX943);
  not NOT_183(WX570,WX945);
  not NOT_184(WX571,WX947);
  not NOT_185(WX572,WX949);
  not NOT_186(WX573,WX951);
  not NOT_187(WX574,WX953);
  not NOT_188(WX575,WX955);
  not NOT_189(WX576,WX957);
  not NOT_190(WX577,WX959);
  not NOT_191(WX578,WX961);
  not NOT_192(WX579,WX963);
  not NOT_193(WX580,WX548);
  not NOT_194(WX581,WX549);
  not NOT_195(WX582,WX550);
  not NOT_196(WX583,WX551);
  not NOT_197(WX584,WX552);
  not NOT_198(WX585,WX553);
  not NOT_199(WX586,WX554);
  not NOT_200(WX587,WX555);
  not NOT_201(WX588,WX556);
  not NOT_202(WX589,WX557);
  not NOT_203(WX590,WX558);
  not NOT_204(WX591,WX559);
  not NOT_205(WX592,WX560);
  not NOT_206(WX593,WX561);
  not NOT_207(WX594,WX562);
  not NOT_208(WX595,WX563);
  not NOT_209(WX596,WX564);
  not NOT_210(WX597,WX565);
  not NOT_211(WX598,WX566);
  not NOT_212(WX599,WX567);
  not NOT_213(WX600,WX568);
  not NOT_214(WX601,WX569);
  not NOT_215(WX602,WX570);
  not NOT_216(WX603,WX571);
  not NOT_217(WX604,WX572);
  not NOT_218(WX605,WX573);
  not NOT_219(WX606,WX574);
  not NOT_220(WX607,WX575);
  not NOT_221(WX608,WX576);
  not NOT_222(WX609,WX577);
  not NOT_223(WX610,WX578);
  not NOT_224(WX611,WX579);
  not NOT_225(WX612,WX837);
  not NOT_226(WX613,WX839);
  not NOT_227(WX614,WX841);
  not NOT_228(WX615,WX843);
  not NOT_229(WX616,WX845);
  not NOT_230(WX617,WX847);
  not NOT_231(WX618,WX849);
  not NOT_232(WX619,WX851);
  not NOT_233(WX620,WX853);
  not NOT_234(WX621,WX855);
  not NOT_235(WX622,WX857);
  not NOT_236(WX623,WX859);
  not NOT_237(WX624,WX861);
  not NOT_238(WX625,WX863);
  not NOT_239(WX626,WX865);
  not NOT_240(WX627,WX867);
  not NOT_241(WX628,WX869);
  not NOT_242(WX629,WX871);
  not NOT_243(WX630,WX873);
  not NOT_244(WX631,WX875);
  not NOT_245(WX632,WX877);
  not NOT_246(WX633,WX879);
  not NOT_247(WX634,WX881);
  not NOT_248(WX635,WX883);
  not NOT_249(WX636,WX885);
  not NOT_250(WX637,WX887);
  not NOT_251(WX638,WX889);
  not NOT_252(WX639,WX891);
  not NOT_253(WX640,WX893);
  not NOT_254(WX641,WX895);
  not NOT_255(WX642,WX897);
  not NOT_256(WX643,WX899);
  not NOT_257(WX932,WX916);
  not NOT_258(WX933,WX932);
  not NOT_259(WX934,WX917);
  not NOT_260(WX935,WX934);
  not NOT_261(WX936,WX918);
  not NOT_262(WX937,WX936);
  not NOT_263(WX938,WX919);
  not NOT_264(WX939,WX938);
  not NOT_265(WX940,WX920);
  not NOT_266(WX941,WX940);
  not NOT_267(WX942,WX921);
  not NOT_268(WX943,WX942);
  not NOT_269(WX944,WX922);
  not NOT_270(WX945,WX944);
  not NOT_271(WX946,WX923);
  not NOT_272(WX947,WX946);
  not NOT_273(WX948,WX924);
  not NOT_274(WX949,WX948);
  not NOT_275(WX950,WX925);
  not NOT_276(WX951,WX950);
  not NOT_277(WX952,WX926);
  not NOT_278(WX953,WX952);
  not NOT_279(WX954,WX927);
  not NOT_280(WX955,WX954);
  not NOT_281(WX956,WX928);
  not NOT_282(WX957,WX956);
  not NOT_283(WX958,WX929);
  not NOT_284(WX959,WX958);
  not NOT_285(WX960,WX930);
  not NOT_286(WX961,WX960);
  not NOT_287(WX962,WX931);
  not NOT_288(WX963,WX962);
  not NOT_289(WX964,WX900);
  not NOT_290(WX965,WX964);
  not NOT_291(WX966,WX901);
  not NOT_292(WX967,WX966);
  not NOT_293(WX968,WX902);
  not NOT_294(WX969,WX968);
  not NOT_295(WX970,WX903);
  not NOT_296(WX971,WX970);
  not NOT_297(WX972,WX904);
  not NOT_298(WX973,WX972);
  not NOT_299(WX974,WX905);
  not NOT_300(WX975,WX974);
  not NOT_301(WX976,WX906);
  not NOT_302(WX977,WX976);
  not NOT_303(WX978,WX907);
  not NOT_304(WX979,WX978);
  not NOT_305(WX980,WX908);
  not NOT_306(WX981,WX980);
  not NOT_307(WX982,WX909);
  not NOT_308(WX983,WX982);
  not NOT_309(WX984,WX910);
  not NOT_310(WX985,WX984);
  not NOT_311(WX986,WX911);
  not NOT_312(WX987,WX986);
  not NOT_313(WX988,WX912);
  not NOT_314(WX989,WX988);
  not NOT_315(WX990,WX913);
  not NOT_316(WX991,WX990);
  not NOT_317(WX992,WX914);
  not NOT_318(WX993,WX992);
  not NOT_319(WX994,WX915);
  not NOT_320(WX995,WX994);
  not NOT_321(WX996,TM0);
  not NOT_322(WX997,TM0);
  not NOT_323(WX998,TM0);
  not NOT_324(WX999,TM1);
  not NOT_325(WX1000,TM1);
  not NOT_326(WX1001,WX1000);
  not NOT_327(WX1002,WX998);
  not NOT_328(WX1003,WX999);
  not NOT_329(WX1004,WX997);
  not NOT_330(WX1005,WX996);
  not NOT_331(WX1009,WX1005);
  not NOT_332(WX1011,WX1010);
  not NOT_333(DATA_9_31,WX1011);
  not NOT_334(WX1016,WX1005);
  not NOT_335(WX1018,WX1017);
  not NOT_336(DATA_9_30,WX1018);
  not NOT_337(WX1023,WX1005);
  not NOT_338(WX1025,WX1024);
  not NOT_339(DATA_9_29,WX1025);
  not NOT_340(WX1030,WX1005);
  not NOT_341(WX1032,WX1031);
  not NOT_342(DATA_9_28,WX1032);
  not NOT_343(WX1037,WX1005);
  not NOT_344(WX1039,WX1038);
  not NOT_345(DATA_9_27,WX1039);
  not NOT_346(WX1044,WX1005);
  not NOT_347(WX1046,WX1045);
  not NOT_348(DATA_9_26,WX1046);
  not NOT_349(WX1051,WX1005);
  not NOT_350(WX1053,WX1052);
  not NOT_351(DATA_9_25,WX1053);
  not NOT_352(WX1058,WX1005);
  not NOT_353(WX1060,WX1059);
  not NOT_354(DATA_9_24,WX1060);
  not NOT_355(WX1065,WX1005);
  not NOT_356(WX1067,WX1066);
  not NOT_357(DATA_9_23,WX1067);
  not NOT_358(WX1072,WX1005);
  not NOT_359(WX1074,WX1073);
  not NOT_360(DATA_9_22,WX1074);
  not NOT_361(WX1079,WX1005);
  not NOT_362(WX1081,WX1080);
  not NOT_363(DATA_9_21,WX1081);
  not NOT_364(WX1086,WX1005);
  not NOT_365(WX1088,WX1087);
  not NOT_366(DATA_9_20,WX1088);
  not NOT_367(WX1093,WX1005);
  not NOT_368(WX1095,WX1094);
  not NOT_369(DATA_9_19,WX1095);
  not NOT_370(WX1100,WX1005);
  not NOT_371(WX1102,WX1101);
  not NOT_372(DATA_9_18,WX1102);
  not NOT_373(WX1107,WX1005);
  not NOT_374(WX1109,WX1108);
  not NOT_375(DATA_9_17,WX1109);
  not NOT_376(WX1114,WX1005);
  not NOT_377(WX1116,WX1115);
  not NOT_378(DATA_9_16,WX1116);
  not NOT_379(WX1121,WX1005);
  not NOT_380(WX1123,WX1122);
  not NOT_381(DATA_9_15,WX1123);
  not NOT_382(WX1128,WX1005);
  not NOT_383(WX1130,WX1129);
  not NOT_384(DATA_9_14,WX1130);
  not NOT_385(WX1135,WX1005);
  not NOT_386(WX1137,WX1136);
  not NOT_387(DATA_9_13,WX1137);
  not NOT_388(WX1142,WX1005);
  not NOT_389(WX1144,WX1143);
  not NOT_390(DATA_9_12,WX1144);
  not NOT_391(WX1149,WX1005);
  not NOT_392(WX1151,WX1150);
  not NOT_393(DATA_9_11,WX1151);
  not NOT_394(WX1156,WX1005);
  not NOT_395(WX1158,WX1157);
  not NOT_396(DATA_9_10,WX1158);
  not NOT_397(WX1163,WX1005);
  not NOT_398(WX1165,WX1164);
  not NOT_399(DATA_9_9,WX1165);
  not NOT_400(WX1170,WX1005);
  not NOT_401(WX1172,WX1171);
  not NOT_402(DATA_9_8,WX1172);
  not NOT_403(WX1177,WX1005);
  not NOT_404(WX1179,WX1178);
  not NOT_405(DATA_9_7,WX1179);
  not NOT_406(WX1184,WX1005);
  not NOT_407(WX1186,WX1185);
  not NOT_408(DATA_9_6,WX1186);
  not NOT_409(WX1191,WX1005);
  not NOT_410(WX1193,WX1192);
  not NOT_411(DATA_9_5,WX1193);
  not NOT_412(WX1198,WX1005);
  not NOT_413(WX1200,WX1199);
  not NOT_414(DATA_9_4,WX1200);
  not NOT_415(WX1205,WX1005);
  not NOT_416(WX1207,WX1206);
  not NOT_417(DATA_9_3,WX1207);
  not NOT_418(WX1212,WX1005);
  not NOT_419(WX1214,WX1213);
  not NOT_420(DATA_9_2,WX1214);
  not NOT_421(WX1219,WX1005);
  not NOT_422(WX1221,WX1220);
  not NOT_423(DATA_9_1,WX1221);
  not NOT_424(WX1226,WX1005);
  not NOT_425(WX1228,WX1227);
  not NOT_426(DATA_9_0,WX1228);
  not NOT_427(WX1230,RESET);
  not NOT_428(WX1263,WX1230);
  not NOT_429(WX1330,WX2296);
  not NOT_430(WX1334,WX2297);
  not NOT_431(WX1338,WX2297);
  not NOT_432(WX1340,WX1331);
  not NOT_433(WX1341,WX1340);
  not NOT_434(WX1344,WX2296);
  not NOT_435(WX1348,WX2297);
  not NOT_436(WX1352,WX2297);
  not NOT_437(WX1354,WX1345);
  not NOT_438(WX1355,WX1354);
  not NOT_439(WX1358,WX2296);
  not NOT_440(WX1362,WX2297);
  not NOT_441(WX1366,WX2297);
  not NOT_442(WX1368,WX1359);
  not NOT_443(WX1369,WX1368);
  not NOT_444(WX1372,WX2296);
  not NOT_445(WX1376,WX2297);
  not NOT_446(WX1380,WX2297);
  not NOT_447(WX1382,WX1373);
  not NOT_448(WX1383,WX1382);
  not NOT_449(WX1386,WX2296);
  not NOT_450(WX1390,WX2297);
  not NOT_451(WX1394,WX2297);
  not NOT_452(WX1396,WX1387);
  not NOT_453(WX1397,WX1396);
  not NOT_454(WX1400,WX2296);
  not NOT_455(WX1404,WX2297);
  not NOT_456(WX1408,WX2297);
  not NOT_457(WX1410,WX1401);
  not NOT_458(WX1411,WX1410);
  not NOT_459(WX1414,WX2296);
  not NOT_460(WX1418,WX2297);
  not NOT_461(WX1422,WX2297);
  not NOT_462(WX1424,WX1415);
  not NOT_463(WX1425,WX1424);
  not NOT_464(WX1428,WX2296);
  not NOT_465(WX1432,WX2297);
  not NOT_466(WX1436,WX2297);
  not NOT_467(WX1438,WX1429);
  not NOT_468(WX1439,WX1438);
  not NOT_469(WX1442,WX2296);
  not NOT_470(WX1446,WX2297);
  not NOT_471(WX1450,WX2297);
  not NOT_472(WX1452,WX1443);
  not NOT_473(WX1453,WX1452);
  not NOT_474(WX1456,WX2296);
  not NOT_475(WX1460,WX2297);
  not NOT_476(WX1464,WX2297);
  not NOT_477(WX1466,WX1457);
  not NOT_478(WX1467,WX1466);
  not NOT_479(WX1470,WX2296);
  not NOT_480(WX1474,WX2297);
  not NOT_481(WX1478,WX2297);
  not NOT_482(WX1480,WX1471);
  not NOT_483(WX1481,WX1480);
  not NOT_484(WX1484,WX2296);
  not NOT_485(WX1488,WX2297);
  not NOT_486(WX1492,WX2297);
  not NOT_487(WX1494,WX1485);
  not NOT_488(WX1495,WX1494);
  not NOT_489(WX1498,WX2296);
  not NOT_490(WX1502,WX2297);
  not NOT_491(WX1506,WX2297);
  not NOT_492(WX1508,WX1499);
  not NOT_493(WX1509,WX1508);
  not NOT_494(WX1512,WX2296);
  not NOT_495(WX1516,WX2297);
  not NOT_496(WX1520,WX2297);
  not NOT_497(WX1522,WX1513);
  not NOT_498(WX1523,WX1522);
  not NOT_499(WX1526,WX2296);
  not NOT_500(WX1530,WX2297);
  not NOT_501(WX1534,WX2297);
  not NOT_502(WX1536,WX1527);
  not NOT_503(WX1537,WX1536);
  not NOT_504(WX1540,WX2296);
  not NOT_505(WX1544,WX2297);
  not NOT_506(WX1548,WX2297);
  not NOT_507(WX1550,WX1541);
  not NOT_508(WX1551,WX1550);
  not NOT_509(WX1554,WX2296);
  not NOT_510(WX1558,WX2297);
  not NOT_511(WX1562,WX2297);
  not NOT_512(WX1564,WX1555);
  not NOT_513(WX1565,WX1564);
  not NOT_514(WX1568,WX2296);
  not NOT_515(WX1572,WX2297);
  not NOT_516(WX1576,WX2297);
  not NOT_517(WX1578,WX1569);
  not NOT_518(WX1579,WX1578);
  not NOT_519(WX1582,WX2296);
  not NOT_520(WX1586,WX2297);
  not NOT_521(WX1590,WX2297);
  not NOT_522(WX1592,WX1583);
  not NOT_523(WX1593,WX1592);
  not NOT_524(WX1596,WX2296);
  not NOT_525(WX1600,WX2297);
  not NOT_526(WX1604,WX2297);
  not NOT_527(WX1606,WX1597);
  not NOT_528(WX1607,WX1606);
  not NOT_529(WX1610,WX2296);
  not NOT_530(WX1614,WX2297);
  not NOT_531(WX1618,WX2297);
  not NOT_532(WX1620,WX1611);
  not NOT_533(WX1621,WX1620);
  not NOT_534(WX1624,WX2296);
  not NOT_535(WX1628,WX2297);
  not NOT_536(WX1632,WX2297);
  not NOT_537(WX1634,WX1625);
  not NOT_538(WX1635,WX1634);
  not NOT_539(WX1638,WX2296);
  not NOT_540(WX1642,WX2297);
  not NOT_541(WX1646,WX2297);
  not NOT_542(WX1648,WX1639);
  not NOT_543(WX1649,WX1648);
  not NOT_544(WX1652,WX2296);
  not NOT_545(WX1656,WX2297);
  not NOT_546(WX1660,WX2297);
  not NOT_547(WX1662,WX1653);
  not NOT_548(WX1663,WX1662);
  not NOT_549(WX1666,WX2296);
  not NOT_550(WX1670,WX2297);
  not NOT_551(WX1674,WX2297);
  not NOT_552(WX1676,WX1667);
  not NOT_553(WX1677,WX1676);
  not NOT_554(WX1680,WX2296);
  not NOT_555(WX1684,WX2297);
  not NOT_556(WX1688,WX2297);
  not NOT_557(WX1690,WX1681);
  not NOT_558(WX1691,WX1690);
  not NOT_559(WX1694,WX2296);
  not NOT_560(WX1698,WX2297);
  not NOT_561(WX1702,WX2297);
  not NOT_562(WX1704,WX1695);
  not NOT_563(WX1705,WX1704);
  not NOT_564(WX1708,WX2296);
  not NOT_565(WX1712,WX2297);
  not NOT_566(WX1716,WX2297);
  not NOT_567(WX1718,WX1709);
  not NOT_568(WX1719,WX1718);
  not NOT_569(WX1722,WX2296);
  not NOT_570(WX1726,WX2297);
  not NOT_571(WX1730,WX2297);
  not NOT_572(WX1732,WX1723);
  not NOT_573(WX1733,WX1732);
  not NOT_574(WX1736,WX2296);
  not NOT_575(WX1740,WX2297);
  not NOT_576(WX1744,WX2297);
  not NOT_577(WX1746,WX1737);
  not NOT_578(WX1747,WX1746);
  not NOT_579(WX1750,WX2296);
  not NOT_580(WX1754,WX2297);
  not NOT_581(WX1758,WX2297);
  not NOT_582(WX1760,WX1751);
  not NOT_583(WX1761,WX1760);
  not NOT_584(WX1764,WX2296);
  not NOT_585(WX1768,WX2297);
  not NOT_586(WX1772,WX2297);
  not NOT_587(WX1774,WX1765);
  not NOT_588(WX1775,WX1774);
  not NOT_589(WX1776,WX1778);
  not NOT_590(WX1841,WX2258);
  not NOT_591(WX1842,WX2260);
  not NOT_592(WX1843,WX2262);
  not NOT_593(WX1844,WX2264);
  not NOT_594(WX1845,WX2266);
  not NOT_595(WX1846,WX2268);
  not NOT_596(WX1847,WX2270);
  not NOT_597(WX1848,WX2272);
  not NOT_598(WX1849,WX2274);
  not NOT_599(WX1850,WX2276);
  not NOT_600(WX1851,WX2278);
  not NOT_601(WX1852,WX2280);
  not NOT_602(WX1853,WX2282);
  not NOT_603(WX1854,WX2284);
  not NOT_604(WX1855,WX2286);
  not NOT_605(WX1856,WX2288);
  not NOT_606(WX1857,WX2226);
  not NOT_607(WX1858,WX2228);
  not NOT_608(WX1859,WX2230);
  not NOT_609(WX1860,WX2232);
  not NOT_610(WX1861,WX2234);
  not NOT_611(WX1862,WX2236);
  not NOT_612(WX1863,WX2238);
  not NOT_613(WX1864,WX2240);
  not NOT_614(WX1865,WX2242);
  not NOT_615(WX1866,WX2244);
  not NOT_616(WX1867,WX2246);
  not NOT_617(WX1868,WX2248);
  not NOT_618(WX1869,WX2250);
  not NOT_619(WX1870,WX2252);
  not NOT_620(WX1871,WX2254);
  not NOT_621(WX1872,WX2256);
  not NOT_622(WX1873,WX1841);
  not NOT_623(WX1874,WX1842);
  not NOT_624(WX1875,WX1843);
  not NOT_625(WX1876,WX1844);
  not NOT_626(WX1877,WX1845);
  not NOT_627(WX1878,WX1846);
  not NOT_628(WX1879,WX1847);
  not NOT_629(WX1880,WX1848);
  not NOT_630(WX1881,WX1849);
  not NOT_631(WX1882,WX1850);
  not NOT_632(WX1883,WX1851);
  not NOT_633(WX1884,WX1852);
  not NOT_634(WX1885,WX1853);
  not NOT_635(WX1886,WX1854);
  not NOT_636(WX1887,WX1855);
  not NOT_637(WX1888,WX1856);
  not NOT_638(WX1889,WX1857);
  not NOT_639(WX1890,WX1858);
  not NOT_640(WX1891,WX1859);
  not NOT_641(WX1892,WX1860);
  not NOT_642(WX1893,WX1861);
  not NOT_643(WX1894,WX1862);
  not NOT_644(WX1895,WX1863);
  not NOT_645(WX1896,WX1864);
  not NOT_646(WX1897,WX1865);
  not NOT_647(WX1898,WX1866);
  not NOT_648(WX1899,WX1867);
  not NOT_649(WX1900,WX1868);
  not NOT_650(WX1901,WX1869);
  not NOT_651(WX1902,WX1870);
  not NOT_652(WX1903,WX1871);
  not NOT_653(WX1904,WX1872);
  not NOT_654(WX1905,WX2130);
  not NOT_655(WX1906,WX2132);
  not NOT_656(WX1907,WX2134);
  not NOT_657(WX1908,WX2136);
  not NOT_658(WX1909,WX2138);
  not NOT_659(WX1910,WX2140);
  not NOT_660(WX1911,WX2142);
  not NOT_661(WX1912,WX2144);
  not NOT_662(WX1913,WX2146);
  not NOT_663(WX1914,WX2148);
  not NOT_664(WX1915,WX2150);
  not NOT_665(WX1916,WX2152);
  not NOT_666(WX1917,WX2154);
  not NOT_667(WX1918,WX2156);
  not NOT_668(WX1919,WX2158);
  not NOT_669(WX1920,WX2160);
  not NOT_670(WX1921,WX2162);
  not NOT_671(WX1922,WX2164);
  not NOT_672(WX1923,WX2166);
  not NOT_673(WX1924,WX2168);
  not NOT_674(WX1925,WX2170);
  not NOT_675(WX1926,WX2172);
  not NOT_676(WX1927,WX2174);
  not NOT_677(WX1928,WX2176);
  not NOT_678(WX1929,WX2178);
  not NOT_679(WX1930,WX2180);
  not NOT_680(WX1931,WX2182);
  not NOT_681(WX1932,WX2184);
  not NOT_682(WX1933,WX2186);
  not NOT_683(WX1934,WX2188);
  not NOT_684(WX1935,WX2190);
  not NOT_685(WX1936,WX2192);
  not NOT_686(WX2225,WX2209);
  not NOT_687(WX2226,WX2225);
  not NOT_688(WX2227,WX2210);
  not NOT_689(WX2228,WX2227);
  not NOT_690(WX2229,WX2211);
  not NOT_691(WX2230,WX2229);
  not NOT_692(WX2231,WX2212);
  not NOT_693(WX2232,WX2231);
  not NOT_694(WX2233,WX2213);
  not NOT_695(WX2234,WX2233);
  not NOT_696(WX2235,WX2214);
  not NOT_697(WX2236,WX2235);
  not NOT_698(WX2237,WX2215);
  not NOT_699(WX2238,WX2237);
  not NOT_700(WX2239,WX2216);
  not NOT_701(WX2240,WX2239);
  not NOT_702(WX2241,WX2217);
  not NOT_703(WX2242,WX2241);
  not NOT_704(WX2243,WX2218);
  not NOT_705(WX2244,WX2243);
  not NOT_706(WX2245,WX2219);
  not NOT_707(WX2246,WX2245);
  not NOT_708(WX2247,WX2220);
  not NOT_709(WX2248,WX2247);
  not NOT_710(WX2249,WX2221);
  not NOT_711(WX2250,WX2249);
  not NOT_712(WX2251,WX2222);
  not NOT_713(WX2252,WX2251);
  not NOT_714(WX2253,WX2223);
  not NOT_715(WX2254,WX2253);
  not NOT_716(WX2255,WX2224);
  not NOT_717(WX2256,WX2255);
  not NOT_718(WX2257,WX2193);
  not NOT_719(WX2258,WX2257);
  not NOT_720(WX2259,WX2194);
  not NOT_721(WX2260,WX2259);
  not NOT_722(WX2261,WX2195);
  not NOT_723(WX2262,WX2261);
  not NOT_724(WX2263,WX2196);
  not NOT_725(WX2264,WX2263);
  not NOT_726(WX2265,WX2197);
  not NOT_727(WX2266,WX2265);
  not NOT_728(WX2267,WX2198);
  not NOT_729(WX2268,WX2267);
  not NOT_730(WX2269,WX2199);
  not NOT_731(WX2270,WX2269);
  not NOT_732(WX2271,WX2200);
  not NOT_733(WX2272,WX2271);
  not NOT_734(WX2273,WX2201);
  not NOT_735(WX2274,WX2273);
  not NOT_736(WX2275,WX2202);
  not NOT_737(WX2276,WX2275);
  not NOT_738(WX2277,WX2203);
  not NOT_739(WX2278,WX2277);
  not NOT_740(WX2279,WX2204);
  not NOT_741(WX2280,WX2279);
  not NOT_742(WX2281,WX2205);
  not NOT_743(WX2282,WX2281);
  not NOT_744(WX2283,WX2206);
  not NOT_745(WX2284,WX2283);
  not NOT_746(WX2285,WX2207);
  not NOT_747(WX2286,WX2285);
  not NOT_748(WX2287,WX2208);
  not NOT_749(WX2288,WX2287);
  not NOT_750(WX2289,TM0);
  not NOT_751(WX2290,TM0);
  not NOT_752(WX2291,TM0);
  not NOT_753(WX2292,TM1);
  not NOT_754(WX2293,TM1);
  not NOT_755(WX2294,WX2293);
  not NOT_756(WX2295,WX2291);
  not NOT_757(WX2296,WX2292);
  not NOT_758(WX2297,WX2290);
  not NOT_759(WX2298,WX2289);
  not NOT_760(WX2302,WX2298);
  not NOT_761(WX2304,WX2303);
  not NOT_762(WX2305,WX2304);
  not NOT_763(WX2309,WX2298);
  not NOT_764(WX2311,WX2310);
  not NOT_765(WX2312,WX2311);
  not NOT_766(WX2316,WX2298);
  not NOT_767(WX2318,WX2317);
  not NOT_768(WX2319,WX2318);
  not NOT_769(WX2323,WX2298);
  not NOT_770(WX2325,WX2324);
  not NOT_771(WX2326,WX2325);
  not NOT_772(WX2330,WX2298);
  not NOT_773(WX2332,WX2331);
  not NOT_774(WX2333,WX2332);
  not NOT_775(WX2337,WX2298);
  not NOT_776(WX2339,WX2338);
  not NOT_777(WX2340,WX2339);
  not NOT_778(WX2344,WX2298);
  not NOT_779(WX2346,WX2345);
  not NOT_780(WX2347,WX2346);
  not NOT_781(WX2351,WX2298);
  not NOT_782(WX2353,WX2352);
  not NOT_783(WX2354,WX2353);
  not NOT_784(WX2358,WX2298);
  not NOT_785(WX2360,WX2359);
  not NOT_786(WX2361,WX2360);
  not NOT_787(WX2365,WX2298);
  not NOT_788(WX2367,WX2366);
  not NOT_789(WX2368,WX2367);
  not NOT_790(WX2372,WX2298);
  not NOT_791(WX2374,WX2373);
  not NOT_792(WX2375,WX2374);
  not NOT_793(WX2379,WX2298);
  not NOT_794(WX2381,WX2380);
  not NOT_795(WX2382,WX2381);
  not NOT_796(WX2386,WX2298);
  not NOT_797(WX2388,WX2387);
  not NOT_798(WX2389,WX2388);
  not NOT_799(WX2393,WX2298);
  not NOT_800(WX2395,WX2394);
  not NOT_801(WX2396,WX2395);
  not NOT_802(WX2400,WX2298);
  not NOT_803(WX2402,WX2401);
  not NOT_804(WX2403,WX2402);
  not NOT_805(WX2407,WX2298);
  not NOT_806(WX2409,WX2408);
  not NOT_807(WX2410,WX2409);
  not NOT_808(WX2414,WX2298);
  not NOT_809(WX2416,WX2415);
  not NOT_810(WX2417,WX2416);
  not NOT_811(WX2421,WX2298);
  not NOT_812(WX2423,WX2422);
  not NOT_813(WX2424,WX2423);
  not NOT_814(WX2428,WX2298);
  not NOT_815(WX2430,WX2429);
  not NOT_816(WX2431,WX2430);
  not NOT_817(WX2435,WX2298);
  not NOT_818(WX2437,WX2436);
  not NOT_819(WX2438,WX2437);
  not NOT_820(WX2442,WX2298);
  not NOT_821(WX2444,WX2443);
  not NOT_822(WX2445,WX2444);
  not NOT_823(WX2449,WX2298);
  not NOT_824(WX2451,WX2450);
  not NOT_825(WX2452,WX2451);
  not NOT_826(WX2456,WX2298);
  not NOT_827(WX2458,WX2457);
  not NOT_828(WX2459,WX2458);
  not NOT_829(WX2463,WX2298);
  not NOT_830(WX2465,WX2464);
  not NOT_831(WX2466,WX2465);
  not NOT_832(WX2470,WX2298);
  not NOT_833(WX2472,WX2471);
  not NOT_834(WX2473,WX2472);
  not NOT_835(WX2477,WX2298);
  not NOT_836(WX2479,WX2478);
  not NOT_837(WX2480,WX2479);
  not NOT_838(WX2484,WX2298);
  not NOT_839(WX2486,WX2485);
  not NOT_840(WX2487,WX2486);
  not NOT_841(WX2491,WX2298);
  not NOT_842(WX2493,WX2492);
  not NOT_843(WX2494,WX2493);
  not NOT_844(WX2498,WX2298);
  not NOT_845(WX2500,WX2499);
  not NOT_846(WX2501,WX2500);
  not NOT_847(WX2505,WX2298);
  not NOT_848(WX2507,WX2506);
  not NOT_849(WX2508,WX2507);
  not NOT_850(WX2512,WX2298);
  not NOT_851(WX2514,WX2513);
  not NOT_852(WX2515,WX2514);
  not NOT_853(WX2519,WX2298);
  not NOT_854(WX2521,WX2520);
  not NOT_855(WX2522,WX2521);
  not NOT_856(WX2523,RESET);
  not NOT_857(WX2556,WX2523);
  not NOT_858(WX2623,WX3589);
  not NOT_859(WX2627,WX3590);
  not NOT_860(WX2631,WX3590);
  not NOT_861(WX2633,WX2624);
  not NOT_862(WX2634,WX2633);
  not NOT_863(WX2637,WX3589);
  not NOT_864(WX2641,WX3590);
  not NOT_865(WX2645,WX3590);
  not NOT_866(WX2647,WX2638);
  not NOT_867(WX2648,WX2647);
  not NOT_868(WX2651,WX3589);
  not NOT_869(WX2655,WX3590);
  not NOT_870(WX2659,WX3590);
  not NOT_871(WX2661,WX2652);
  not NOT_872(WX2662,WX2661);
  not NOT_873(WX2665,WX3589);
  not NOT_874(WX2669,WX3590);
  not NOT_875(WX2673,WX3590);
  not NOT_876(WX2675,WX2666);
  not NOT_877(WX2676,WX2675);
  not NOT_878(WX2679,WX3589);
  not NOT_879(WX2683,WX3590);
  not NOT_880(WX2687,WX3590);
  not NOT_881(WX2689,WX2680);
  not NOT_882(WX2690,WX2689);
  not NOT_883(WX2693,WX3589);
  not NOT_884(WX2697,WX3590);
  not NOT_885(WX2701,WX3590);
  not NOT_886(WX2703,WX2694);
  not NOT_887(WX2704,WX2703);
  not NOT_888(WX2707,WX3589);
  not NOT_889(WX2711,WX3590);
  not NOT_890(WX2715,WX3590);
  not NOT_891(WX2717,WX2708);
  not NOT_892(WX2718,WX2717);
  not NOT_893(WX2721,WX3589);
  not NOT_894(WX2725,WX3590);
  not NOT_895(WX2729,WX3590);
  not NOT_896(WX2731,WX2722);
  not NOT_897(WX2732,WX2731);
  not NOT_898(WX2735,WX3589);
  not NOT_899(WX2739,WX3590);
  not NOT_900(WX2743,WX3590);
  not NOT_901(WX2745,WX2736);
  not NOT_902(WX2746,WX2745);
  not NOT_903(WX2749,WX3589);
  not NOT_904(WX2753,WX3590);
  not NOT_905(WX2757,WX3590);
  not NOT_906(WX2759,WX2750);
  not NOT_907(WX2760,WX2759);
  not NOT_908(WX2763,WX3589);
  not NOT_909(WX2767,WX3590);
  not NOT_910(WX2771,WX3590);
  not NOT_911(WX2773,WX2764);
  not NOT_912(WX2774,WX2773);
  not NOT_913(WX2777,WX3589);
  not NOT_914(WX2781,WX3590);
  not NOT_915(WX2785,WX3590);
  not NOT_916(WX2787,WX2778);
  not NOT_917(WX2788,WX2787);
  not NOT_918(WX2791,WX3589);
  not NOT_919(WX2795,WX3590);
  not NOT_920(WX2799,WX3590);
  not NOT_921(WX2801,WX2792);
  not NOT_922(WX2802,WX2801);
  not NOT_923(WX2805,WX3589);
  not NOT_924(WX2809,WX3590);
  not NOT_925(WX2813,WX3590);
  not NOT_926(WX2815,WX2806);
  not NOT_927(WX2816,WX2815);
  not NOT_928(WX2819,WX3589);
  not NOT_929(WX2823,WX3590);
  not NOT_930(WX2827,WX3590);
  not NOT_931(WX2829,WX2820);
  not NOT_932(WX2830,WX2829);
  not NOT_933(WX2833,WX3589);
  not NOT_934(WX2837,WX3590);
  not NOT_935(WX2841,WX3590);
  not NOT_936(WX2843,WX2834);
  not NOT_937(WX2844,WX2843);
  not NOT_938(WX2847,WX3589);
  not NOT_939(WX2851,WX3590);
  not NOT_940(WX2855,WX3590);
  not NOT_941(WX2857,WX2848);
  not NOT_942(WX2858,WX2857);
  not NOT_943(WX2861,WX3589);
  not NOT_944(WX2865,WX3590);
  not NOT_945(WX2869,WX3590);
  not NOT_946(WX2871,WX2862);
  not NOT_947(WX2872,WX2871);
  not NOT_948(WX2875,WX3589);
  not NOT_949(WX2879,WX3590);
  not NOT_950(WX2883,WX3590);
  not NOT_951(WX2885,WX2876);
  not NOT_952(WX2886,WX2885);
  not NOT_953(WX2889,WX3589);
  not NOT_954(WX2893,WX3590);
  not NOT_955(WX2897,WX3590);
  not NOT_956(WX2899,WX2890);
  not NOT_957(WX2900,WX2899);
  not NOT_958(WX2903,WX3589);
  not NOT_959(WX2907,WX3590);
  not NOT_960(WX2911,WX3590);
  not NOT_961(WX2913,WX2904);
  not NOT_962(WX2914,WX2913);
  not NOT_963(WX2917,WX3589);
  not NOT_964(WX2921,WX3590);
  not NOT_965(WX2925,WX3590);
  not NOT_966(WX2927,WX2918);
  not NOT_967(WX2928,WX2927);
  not NOT_968(WX2931,WX3589);
  not NOT_969(WX2935,WX3590);
  not NOT_970(WX2939,WX3590);
  not NOT_971(WX2941,WX2932);
  not NOT_972(WX2942,WX2941);
  not NOT_973(WX2945,WX3589);
  not NOT_974(WX2949,WX3590);
  not NOT_975(WX2953,WX3590);
  not NOT_976(WX2955,WX2946);
  not NOT_977(WX2956,WX2955);
  not NOT_978(WX2959,WX3589);
  not NOT_979(WX2963,WX3590);
  not NOT_980(WX2967,WX3590);
  not NOT_981(WX2969,WX2960);
  not NOT_982(WX2970,WX2969);
  not NOT_983(WX2973,WX3589);
  not NOT_984(WX2977,WX3590);
  not NOT_985(WX2981,WX3590);
  not NOT_986(WX2983,WX2974);
  not NOT_987(WX2984,WX2983);
  not NOT_988(WX2987,WX3589);
  not NOT_989(WX2991,WX3590);
  not NOT_990(WX2995,WX3590);
  not NOT_991(WX2997,WX2988);
  not NOT_992(WX2998,WX2997);
  not NOT_993(WX3001,WX3589);
  not NOT_994(WX3005,WX3590);
  not NOT_995(WX3009,WX3590);
  not NOT_996(WX3011,WX3002);
  not NOT_997(WX3012,WX3011);
  not NOT_998(WX3015,WX3589);
  not NOT_999(WX3019,WX3590);
  not NOT_1000(WX3023,WX3590);
  not NOT_1001(WX3025,WX3016);
  not NOT_1002(WX3026,WX3025);
  not NOT_1003(WX3029,WX3589);
  not NOT_1004(WX3033,WX3590);
  not NOT_1005(WX3037,WX3590);
  not NOT_1006(WX3039,WX3030);
  not NOT_1007(WX3040,WX3039);
  not NOT_1008(WX3043,WX3589);
  not NOT_1009(WX3047,WX3590);
  not NOT_1010(WX3051,WX3590);
  not NOT_1011(WX3053,WX3044);
  not NOT_1012(WX3054,WX3053);
  not NOT_1013(WX3057,WX3589);
  not NOT_1014(WX3061,WX3590);
  not NOT_1015(WX3065,WX3590);
  not NOT_1016(WX3067,WX3058);
  not NOT_1017(WX3068,WX3067);
  not NOT_1018(WX3069,WX3071);
  not NOT_1019(WX3134,WX3551);
  not NOT_1020(WX3135,WX3553);
  not NOT_1021(WX3136,WX3555);
  not NOT_1022(WX3137,WX3557);
  not NOT_1023(WX3138,WX3559);
  not NOT_1024(WX3139,WX3561);
  not NOT_1025(WX3140,WX3563);
  not NOT_1026(WX3141,WX3565);
  not NOT_1027(WX3142,WX3567);
  not NOT_1028(WX3143,WX3569);
  not NOT_1029(WX3144,WX3571);
  not NOT_1030(WX3145,WX3573);
  not NOT_1031(WX3146,WX3575);
  not NOT_1032(WX3147,WX3577);
  not NOT_1033(WX3148,WX3579);
  not NOT_1034(WX3149,WX3581);
  not NOT_1035(WX3150,WX3519);
  not NOT_1036(WX3151,WX3521);
  not NOT_1037(WX3152,WX3523);
  not NOT_1038(WX3153,WX3525);
  not NOT_1039(WX3154,WX3527);
  not NOT_1040(WX3155,WX3529);
  not NOT_1041(WX3156,WX3531);
  not NOT_1042(WX3157,WX3533);
  not NOT_1043(WX3158,WX3535);
  not NOT_1044(WX3159,WX3537);
  not NOT_1045(WX3160,WX3539);
  not NOT_1046(WX3161,WX3541);
  not NOT_1047(WX3162,WX3543);
  not NOT_1048(WX3163,WX3545);
  not NOT_1049(WX3164,WX3547);
  not NOT_1050(WX3165,WX3549);
  not NOT_1051(WX3166,WX3134);
  not NOT_1052(WX3167,WX3135);
  not NOT_1053(WX3168,WX3136);
  not NOT_1054(WX3169,WX3137);
  not NOT_1055(WX3170,WX3138);
  not NOT_1056(WX3171,WX3139);
  not NOT_1057(WX3172,WX3140);
  not NOT_1058(WX3173,WX3141);
  not NOT_1059(WX3174,WX3142);
  not NOT_1060(WX3175,WX3143);
  not NOT_1061(WX3176,WX3144);
  not NOT_1062(WX3177,WX3145);
  not NOT_1063(WX3178,WX3146);
  not NOT_1064(WX3179,WX3147);
  not NOT_1065(WX3180,WX3148);
  not NOT_1066(WX3181,WX3149);
  not NOT_1067(WX3182,WX3150);
  not NOT_1068(WX3183,WX3151);
  not NOT_1069(WX3184,WX3152);
  not NOT_1070(WX3185,WX3153);
  not NOT_1071(WX3186,WX3154);
  not NOT_1072(WX3187,WX3155);
  not NOT_1073(WX3188,WX3156);
  not NOT_1074(WX3189,WX3157);
  not NOT_1075(WX3190,WX3158);
  not NOT_1076(WX3191,WX3159);
  not NOT_1077(WX3192,WX3160);
  not NOT_1078(WX3193,WX3161);
  not NOT_1079(WX3194,WX3162);
  not NOT_1080(WX3195,WX3163);
  not NOT_1081(WX3196,WX3164);
  not NOT_1082(WX3197,WX3165);
  not NOT_1083(WX3198,WX3423);
  not NOT_1084(WX3199,WX3425);
  not NOT_1085(WX3200,WX3427);
  not NOT_1086(WX3201,WX3429);
  not NOT_1087(WX3202,WX3431);
  not NOT_1088(WX3203,WX3433);
  not NOT_1089(WX3204,WX3435);
  not NOT_1090(WX3205,WX3437);
  not NOT_1091(WX3206,WX3439);
  not NOT_1092(WX3207,WX3441);
  not NOT_1093(WX3208,WX3443);
  not NOT_1094(WX3209,WX3445);
  not NOT_1095(WX3210,WX3447);
  not NOT_1096(WX3211,WX3449);
  not NOT_1097(WX3212,WX3451);
  not NOT_1098(WX3213,WX3453);
  not NOT_1099(WX3214,WX3455);
  not NOT_1100(WX3215,WX3457);
  not NOT_1101(WX3216,WX3459);
  not NOT_1102(WX3217,WX3461);
  not NOT_1103(WX3218,WX3463);
  not NOT_1104(WX3219,WX3465);
  not NOT_1105(WX3220,WX3467);
  not NOT_1106(WX3221,WX3469);
  not NOT_1107(WX3222,WX3471);
  not NOT_1108(WX3223,WX3473);
  not NOT_1109(WX3224,WX3475);
  not NOT_1110(WX3225,WX3477);
  not NOT_1111(WX3226,WX3479);
  not NOT_1112(WX3227,WX3481);
  not NOT_1113(WX3228,WX3483);
  not NOT_1114(WX3229,WX3485);
  not NOT_1115(WX3518,WX3502);
  not NOT_1116(WX3519,WX3518);
  not NOT_1117(WX3520,WX3503);
  not NOT_1118(WX3521,WX3520);
  not NOT_1119(WX3522,WX3504);
  not NOT_1120(WX3523,WX3522);
  not NOT_1121(WX3524,WX3505);
  not NOT_1122(WX3525,WX3524);
  not NOT_1123(WX3526,WX3506);
  not NOT_1124(WX3527,WX3526);
  not NOT_1125(WX3528,WX3507);
  not NOT_1126(WX3529,WX3528);
  not NOT_1127(WX3530,WX3508);
  not NOT_1128(WX3531,WX3530);
  not NOT_1129(WX3532,WX3509);
  not NOT_1130(WX3533,WX3532);
  not NOT_1131(WX3534,WX3510);
  not NOT_1132(WX3535,WX3534);
  not NOT_1133(WX3536,WX3511);
  not NOT_1134(WX3537,WX3536);
  not NOT_1135(WX3538,WX3512);
  not NOT_1136(WX3539,WX3538);
  not NOT_1137(WX3540,WX3513);
  not NOT_1138(WX3541,WX3540);
  not NOT_1139(WX3542,WX3514);
  not NOT_1140(WX3543,WX3542);
  not NOT_1141(WX3544,WX3515);
  not NOT_1142(WX3545,WX3544);
  not NOT_1143(WX3546,WX3516);
  not NOT_1144(WX3547,WX3546);
  not NOT_1145(WX3548,WX3517);
  not NOT_1146(WX3549,WX3548);
  not NOT_1147(WX3550,WX3486);
  not NOT_1148(WX3551,WX3550);
  not NOT_1149(WX3552,WX3487);
  not NOT_1150(WX3553,WX3552);
  not NOT_1151(WX3554,WX3488);
  not NOT_1152(WX3555,WX3554);
  not NOT_1153(WX3556,WX3489);
  not NOT_1154(WX3557,WX3556);
  not NOT_1155(WX3558,WX3490);
  not NOT_1156(WX3559,WX3558);
  not NOT_1157(WX3560,WX3491);
  not NOT_1158(WX3561,WX3560);
  not NOT_1159(WX3562,WX3492);
  not NOT_1160(WX3563,WX3562);
  not NOT_1161(WX3564,WX3493);
  not NOT_1162(WX3565,WX3564);
  not NOT_1163(WX3566,WX3494);
  not NOT_1164(WX3567,WX3566);
  not NOT_1165(WX3568,WX3495);
  not NOT_1166(WX3569,WX3568);
  not NOT_1167(WX3570,WX3496);
  not NOT_1168(WX3571,WX3570);
  not NOT_1169(WX3572,WX3497);
  not NOT_1170(WX3573,WX3572);
  not NOT_1171(WX3574,WX3498);
  not NOT_1172(WX3575,WX3574);
  not NOT_1173(WX3576,WX3499);
  not NOT_1174(WX3577,WX3576);
  not NOT_1175(WX3578,WX3500);
  not NOT_1176(WX3579,WX3578);
  not NOT_1177(WX3580,WX3501);
  not NOT_1178(WX3581,WX3580);
  not NOT_1179(WX3582,TM0);
  not NOT_1180(WX3583,TM0);
  not NOT_1181(WX3584,TM0);
  not NOT_1182(WX3585,TM1);
  not NOT_1183(WX3586,TM1);
  not NOT_1184(WX3587,WX3586);
  not NOT_1185(WX3588,WX3584);
  not NOT_1186(WX3589,WX3585);
  not NOT_1187(WX3590,WX3583);
  not NOT_1188(WX3591,WX3582);
  not NOT_1189(WX3595,WX3591);
  not NOT_1190(WX3597,WX3596);
  not NOT_1191(WX3598,WX3597);
  not NOT_1192(WX3602,WX3591);
  not NOT_1193(WX3604,WX3603);
  not NOT_1194(WX3605,WX3604);
  not NOT_1195(WX3609,WX3591);
  not NOT_1196(WX3611,WX3610);
  not NOT_1197(WX3612,WX3611);
  not NOT_1198(WX3616,WX3591);
  not NOT_1199(WX3618,WX3617);
  not NOT_1200(WX3619,WX3618);
  not NOT_1201(WX3623,WX3591);
  not NOT_1202(WX3625,WX3624);
  not NOT_1203(WX3626,WX3625);
  not NOT_1204(WX3630,WX3591);
  not NOT_1205(WX3632,WX3631);
  not NOT_1206(WX3633,WX3632);
  not NOT_1207(WX3637,WX3591);
  not NOT_1208(WX3639,WX3638);
  not NOT_1209(WX3640,WX3639);
  not NOT_1210(WX3644,WX3591);
  not NOT_1211(WX3646,WX3645);
  not NOT_1212(WX3647,WX3646);
  not NOT_1213(WX3651,WX3591);
  not NOT_1214(WX3653,WX3652);
  not NOT_1215(WX3654,WX3653);
  not NOT_1216(WX3658,WX3591);
  not NOT_1217(WX3660,WX3659);
  not NOT_1218(WX3661,WX3660);
  not NOT_1219(WX3665,WX3591);
  not NOT_1220(WX3667,WX3666);
  not NOT_1221(WX3668,WX3667);
  not NOT_1222(WX3672,WX3591);
  not NOT_1223(WX3674,WX3673);
  not NOT_1224(WX3675,WX3674);
  not NOT_1225(WX3679,WX3591);
  not NOT_1226(WX3681,WX3680);
  not NOT_1227(WX3682,WX3681);
  not NOT_1228(WX3686,WX3591);
  not NOT_1229(WX3688,WX3687);
  not NOT_1230(WX3689,WX3688);
  not NOT_1231(WX3693,WX3591);
  not NOT_1232(WX3695,WX3694);
  not NOT_1233(WX3696,WX3695);
  not NOT_1234(WX3700,WX3591);
  not NOT_1235(WX3702,WX3701);
  not NOT_1236(WX3703,WX3702);
  not NOT_1237(WX3707,WX3591);
  not NOT_1238(WX3709,WX3708);
  not NOT_1239(WX3710,WX3709);
  not NOT_1240(WX3714,WX3591);
  not NOT_1241(WX3716,WX3715);
  not NOT_1242(WX3717,WX3716);
  not NOT_1243(WX3721,WX3591);
  not NOT_1244(WX3723,WX3722);
  not NOT_1245(WX3724,WX3723);
  not NOT_1246(WX3728,WX3591);
  not NOT_1247(WX3730,WX3729);
  not NOT_1248(WX3731,WX3730);
  not NOT_1249(WX3735,WX3591);
  not NOT_1250(WX3737,WX3736);
  not NOT_1251(WX3738,WX3737);
  not NOT_1252(WX3742,WX3591);
  not NOT_1253(WX3744,WX3743);
  not NOT_1254(WX3745,WX3744);
  not NOT_1255(WX3749,WX3591);
  not NOT_1256(WX3751,WX3750);
  not NOT_1257(WX3752,WX3751);
  not NOT_1258(WX3756,WX3591);
  not NOT_1259(WX3758,WX3757);
  not NOT_1260(WX3759,WX3758);
  not NOT_1261(WX3763,WX3591);
  not NOT_1262(WX3765,WX3764);
  not NOT_1263(WX3766,WX3765);
  not NOT_1264(WX3770,WX3591);
  not NOT_1265(WX3772,WX3771);
  not NOT_1266(WX3773,WX3772);
  not NOT_1267(WX3777,WX3591);
  not NOT_1268(WX3779,WX3778);
  not NOT_1269(WX3780,WX3779);
  not NOT_1270(WX3784,WX3591);
  not NOT_1271(WX3786,WX3785);
  not NOT_1272(WX3787,WX3786);
  not NOT_1273(WX3791,WX3591);
  not NOT_1274(WX3793,WX3792);
  not NOT_1275(WX3794,WX3793);
  not NOT_1276(WX3798,WX3591);
  not NOT_1277(WX3800,WX3799);
  not NOT_1278(WX3801,WX3800);
  not NOT_1279(WX3805,WX3591);
  not NOT_1280(WX3807,WX3806);
  not NOT_1281(WX3808,WX3807);
  not NOT_1282(WX3812,WX3591);
  not NOT_1283(WX3814,WX3813);
  not NOT_1284(WX3815,WX3814);
  not NOT_1285(WX3816,RESET);
  not NOT_1286(WX3849,WX3816);
  not NOT_1287(WX3916,WX4882);
  not NOT_1288(WX3920,WX4883);
  not NOT_1289(WX3924,WX4883);
  not NOT_1290(WX3926,WX3917);
  not NOT_1291(WX3927,WX3926);
  not NOT_1292(WX3930,WX4882);
  not NOT_1293(WX3934,WX4883);
  not NOT_1294(WX3938,WX4883);
  not NOT_1295(WX3940,WX3931);
  not NOT_1296(WX3941,WX3940);
  not NOT_1297(WX3944,WX4882);
  not NOT_1298(WX3948,WX4883);
  not NOT_1299(WX3952,WX4883);
  not NOT_1300(WX3954,WX3945);
  not NOT_1301(WX3955,WX3954);
  not NOT_1302(WX3958,WX4882);
  not NOT_1303(WX3962,WX4883);
  not NOT_1304(WX3966,WX4883);
  not NOT_1305(WX3968,WX3959);
  not NOT_1306(WX3969,WX3968);
  not NOT_1307(WX3972,WX4882);
  not NOT_1308(WX3976,WX4883);
  not NOT_1309(WX3980,WX4883);
  not NOT_1310(WX3982,WX3973);
  not NOT_1311(WX3983,WX3982);
  not NOT_1312(WX3986,WX4882);
  not NOT_1313(WX3990,WX4883);
  not NOT_1314(WX3994,WX4883);
  not NOT_1315(WX3996,WX3987);
  not NOT_1316(WX3997,WX3996);
  not NOT_1317(WX4000,WX4882);
  not NOT_1318(WX4004,WX4883);
  not NOT_1319(WX4008,WX4883);
  not NOT_1320(WX4010,WX4001);
  not NOT_1321(WX4011,WX4010);
  not NOT_1322(WX4014,WX4882);
  not NOT_1323(WX4018,WX4883);
  not NOT_1324(WX4022,WX4883);
  not NOT_1325(WX4024,WX4015);
  not NOT_1326(WX4025,WX4024);
  not NOT_1327(WX4028,WX4882);
  not NOT_1328(WX4032,WX4883);
  not NOT_1329(WX4036,WX4883);
  not NOT_1330(WX4038,WX4029);
  not NOT_1331(WX4039,WX4038);
  not NOT_1332(WX4042,WX4882);
  not NOT_1333(WX4046,WX4883);
  not NOT_1334(WX4050,WX4883);
  not NOT_1335(WX4052,WX4043);
  not NOT_1336(WX4053,WX4052);
  not NOT_1337(WX4056,WX4882);
  not NOT_1338(WX4060,WX4883);
  not NOT_1339(WX4064,WX4883);
  not NOT_1340(WX4066,WX4057);
  not NOT_1341(WX4067,WX4066);
  not NOT_1342(WX4070,WX4882);
  not NOT_1343(WX4074,WX4883);
  not NOT_1344(WX4078,WX4883);
  not NOT_1345(WX4080,WX4071);
  not NOT_1346(WX4081,WX4080);
  not NOT_1347(WX4084,WX4882);
  not NOT_1348(WX4088,WX4883);
  not NOT_1349(WX4092,WX4883);
  not NOT_1350(WX4094,WX4085);
  not NOT_1351(WX4095,WX4094);
  not NOT_1352(WX4098,WX4882);
  not NOT_1353(WX4102,WX4883);
  not NOT_1354(WX4106,WX4883);
  not NOT_1355(WX4108,WX4099);
  not NOT_1356(WX4109,WX4108);
  not NOT_1357(WX4112,WX4882);
  not NOT_1358(WX4116,WX4883);
  not NOT_1359(WX4120,WX4883);
  not NOT_1360(WX4122,WX4113);
  not NOT_1361(WX4123,WX4122);
  not NOT_1362(WX4126,WX4882);
  not NOT_1363(WX4130,WX4883);
  not NOT_1364(WX4134,WX4883);
  not NOT_1365(WX4136,WX4127);
  not NOT_1366(WX4137,WX4136);
  not NOT_1367(WX4140,WX4882);
  not NOT_1368(WX4144,WX4883);
  not NOT_1369(WX4148,WX4883);
  not NOT_1370(WX4150,WX4141);
  not NOT_1371(WX4151,WX4150);
  not NOT_1372(WX4154,WX4882);
  not NOT_1373(WX4158,WX4883);
  not NOT_1374(WX4162,WX4883);
  not NOT_1375(WX4164,WX4155);
  not NOT_1376(WX4165,WX4164);
  not NOT_1377(WX4168,WX4882);
  not NOT_1378(WX4172,WX4883);
  not NOT_1379(WX4176,WX4883);
  not NOT_1380(WX4178,WX4169);
  not NOT_1381(WX4179,WX4178);
  not NOT_1382(WX4182,WX4882);
  not NOT_1383(WX4186,WX4883);
  not NOT_1384(WX4190,WX4883);
  not NOT_1385(WX4192,WX4183);
  not NOT_1386(WX4193,WX4192);
  not NOT_1387(WX4196,WX4882);
  not NOT_1388(WX4200,WX4883);
  not NOT_1389(WX4204,WX4883);
  not NOT_1390(WX4206,WX4197);
  not NOT_1391(WX4207,WX4206);
  not NOT_1392(WX4210,WX4882);
  not NOT_1393(WX4214,WX4883);
  not NOT_1394(WX4218,WX4883);
  not NOT_1395(WX4220,WX4211);
  not NOT_1396(WX4221,WX4220);
  not NOT_1397(WX4224,WX4882);
  not NOT_1398(WX4228,WX4883);
  not NOT_1399(WX4232,WX4883);
  not NOT_1400(WX4234,WX4225);
  not NOT_1401(WX4235,WX4234);
  not NOT_1402(WX4238,WX4882);
  not NOT_1403(WX4242,WX4883);
  not NOT_1404(WX4246,WX4883);
  not NOT_1405(WX4248,WX4239);
  not NOT_1406(WX4249,WX4248);
  not NOT_1407(WX4252,WX4882);
  not NOT_1408(WX4256,WX4883);
  not NOT_1409(WX4260,WX4883);
  not NOT_1410(WX4262,WX4253);
  not NOT_1411(WX4263,WX4262);
  not NOT_1412(WX4266,WX4882);
  not NOT_1413(WX4270,WX4883);
  not NOT_1414(WX4274,WX4883);
  not NOT_1415(WX4276,WX4267);
  not NOT_1416(WX4277,WX4276);
  not NOT_1417(WX4280,WX4882);
  not NOT_1418(WX4284,WX4883);
  not NOT_1419(WX4288,WX4883);
  not NOT_1420(WX4290,WX4281);
  not NOT_1421(WX4291,WX4290);
  not NOT_1422(WX4294,WX4882);
  not NOT_1423(WX4298,WX4883);
  not NOT_1424(WX4302,WX4883);
  not NOT_1425(WX4304,WX4295);
  not NOT_1426(WX4305,WX4304);
  not NOT_1427(WX4308,WX4882);
  not NOT_1428(WX4312,WX4883);
  not NOT_1429(WX4316,WX4883);
  not NOT_1430(WX4318,WX4309);
  not NOT_1431(WX4319,WX4318);
  not NOT_1432(WX4322,WX4882);
  not NOT_1433(WX4326,WX4883);
  not NOT_1434(WX4330,WX4883);
  not NOT_1435(WX4332,WX4323);
  not NOT_1436(WX4333,WX4332);
  not NOT_1437(WX4336,WX4882);
  not NOT_1438(WX4340,WX4883);
  not NOT_1439(WX4344,WX4883);
  not NOT_1440(WX4346,WX4337);
  not NOT_1441(WX4347,WX4346);
  not NOT_1442(WX4350,WX4882);
  not NOT_1443(WX4354,WX4883);
  not NOT_1444(WX4358,WX4883);
  not NOT_1445(WX4360,WX4351);
  not NOT_1446(WX4361,WX4360);
  not NOT_1447(WX4362,WX4364);
  not NOT_1448(WX4427,WX4844);
  not NOT_1449(WX4428,WX4846);
  not NOT_1450(WX4429,WX4848);
  not NOT_1451(WX4430,WX4850);
  not NOT_1452(WX4431,WX4852);
  not NOT_1453(WX4432,WX4854);
  not NOT_1454(WX4433,WX4856);
  not NOT_1455(WX4434,WX4858);
  not NOT_1456(WX4435,WX4860);
  not NOT_1457(WX4436,WX4862);
  not NOT_1458(WX4437,WX4864);
  not NOT_1459(WX4438,WX4866);
  not NOT_1460(WX4439,WX4868);
  not NOT_1461(WX4440,WX4870);
  not NOT_1462(WX4441,WX4872);
  not NOT_1463(WX4442,WX4874);
  not NOT_1464(WX4443,WX4812);
  not NOT_1465(WX4444,WX4814);
  not NOT_1466(WX4445,WX4816);
  not NOT_1467(WX4446,WX4818);
  not NOT_1468(WX4447,WX4820);
  not NOT_1469(WX4448,WX4822);
  not NOT_1470(WX4449,WX4824);
  not NOT_1471(WX4450,WX4826);
  not NOT_1472(WX4451,WX4828);
  not NOT_1473(WX4452,WX4830);
  not NOT_1474(WX4453,WX4832);
  not NOT_1475(WX4454,WX4834);
  not NOT_1476(WX4455,WX4836);
  not NOT_1477(WX4456,WX4838);
  not NOT_1478(WX4457,WX4840);
  not NOT_1479(WX4458,WX4842);
  not NOT_1480(WX4459,WX4427);
  not NOT_1481(WX4460,WX4428);
  not NOT_1482(WX4461,WX4429);
  not NOT_1483(WX4462,WX4430);
  not NOT_1484(WX4463,WX4431);
  not NOT_1485(WX4464,WX4432);
  not NOT_1486(WX4465,WX4433);
  not NOT_1487(WX4466,WX4434);
  not NOT_1488(WX4467,WX4435);
  not NOT_1489(WX4468,WX4436);
  not NOT_1490(WX4469,WX4437);
  not NOT_1491(WX4470,WX4438);
  not NOT_1492(WX4471,WX4439);
  not NOT_1493(WX4472,WX4440);
  not NOT_1494(WX4473,WX4441);
  not NOT_1495(WX4474,WX4442);
  not NOT_1496(WX4475,WX4443);
  not NOT_1497(WX4476,WX4444);
  not NOT_1498(WX4477,WX4445);
  not NOT_1499(WX4478,WX4446);
  not NOT_1500(WX4479,WX4447);
  not NOT_1501(WX4480,WX4448);
  not NOT_1502(WX4481,WX4449);
  not NOT_1503(WX4482,WX4450);
  not NOT_1504(WX4483,WX4451);
  not NOT_1505(WX4484,WX4452);
  not NOT_1506(WX4485,WX4453);
  not NOT_1507(WX4486,WX4454);
  not NOT_1508(WX4487,WX4455);
  not NOT_1509(WX4488,WX4456);
  not NOT_1510(WX4489,WX4457);
  not NOT_1511(WX4490,WX4458);
  not NOT_1512(WX4491,WX4716);
  not NOT_1513(WX4492,WX4718);
  not NOT_1514(WX4493,WX4720);
  not NOT_1515(WX4494,WX4722);
  not NOT_1516(WX4495,WX4724);
  not NOT_1517(WX4496,WX4726);
  not NOT_1518(WX4497,WX4728);
  not NOT_1519(WX4498,WX4730);
  not NOT_1520(WX4499,WX4732);
  not NOT_1521(WX4500,WX4734);
  not NOT_1522(WX4501,WX4736);
  not NOT_1523(WX4502,WX4738);
  not NOT_1524(WX4503,WX4740);
  not NOT_1525(WX4504,WX4742);
  not NOT_1526(WX4505,WX4744);
  not NOT_1527(WX4506,WX4746);
  not NOT_1528(WX4507,WX4748);
  not NOT_1529(WX4508,WX4750);
  not NOT_1530(WX4509,WX4752);
  not NOT_1531(WX4510,WX4754);
  not NOT_1532(WX4511,WX4756);
  not NOT_1533(WX4512,WX4758);
  not NOT_1534(WX4513,WX4760);
  not NOT_1535(WX4514,WX4762);
  not NOT_1536(WX4515,WX4764);
  not NOT_1537(WX4516,WX4766);
  not NOT_1538(WX4517,WX4768);
  not NOT_1539(WX4518,WX4770);
  not NOT_1540(WX4519,WX4772);
  not NOT_1541(WX4520,WX4774);
  not NOT_1542(WX4521,WX4776);
  not NOT_1543(WX4522,WX4778);
  not NOT_1544(WX4811,WX4795);
  not NOT_1545(WX4812,WX4811);
  not NOT_1546(WX4813,WX4796);
  not NOT_1547(WX4814,WX4813);
  not NOT_1548(WX4815,WX4797);
  not NOT_1549(WX4816,WX4815);
  not NOT_1550(WX4817,WX4798);
  not NOT_1551(WX4818,WX4817);
  not NOT_1552(WX4819,WX4799);
  not NOT_1553(WX4820,WX4819);
  not NOT_1554(WX4821,WX4800);
  not NOT_1555(WX4822,WX4821);
  not NOT_1556(WX4823,WX4801);
  not NOT_1557(WX4824,WX4823);
  not NOT_1558(WX4825,WX4802);
  not NOT_1559(WX4826,WX4825);
  not NOT_1560(WX4827,WX4803);
  not NOT_1561(WX4828,WX4827);
  not NOT_1562(WX4829,WX4804);
  not NOT_1563(WX4830,WX4829);
  not NOT_1564(WX4831,WX4805);
  not NOT_1565(WX4832,WX4831);
  not NOT_1566(WX4833,WX4806);
  not NOT_1567(WX4834,WX4833);
  not NOT_1568(WX4835,WX4807);
  not NOT_1569(WX4836,WX4835);
  not NOT_1570(WX4837,WX4808);
  not NOT_1571(WX4838,WX4837);
  not NOT_1572(WX4839,WX4809);
  not NOT_1573(WX4840,WX4839);
  not NOT_1574(WX4841,WX4810);
  not NOT_1575(WX4842,WX4841);
  not NOT_1576(WX4843,WX4779);
  not NOT_1577(WX4844,WX4843);
  not NOT_1578(WX4845,WX4780);
  not NOT_1579(WX4846,WX4845);
  not NOT_1580(WX4847,WX4781);
  not NOT_1581(WX4848,WX4847);
  not NOT_1582(WX4849,WX4782);
  not NOT_1583(WX4850,WX4849);
  not NOT_1584(WX4851,WX4783);
  not NOT_1585(WX4852,WX4851);
  not NOT_1586(WX4853,WX4784);
  not NOT_1587(WX4854,WX4853);
  not NOT_1588(WX4855,WX4785);
  not NOT_1589(WX4856,WX4855);
  not NOT_1590(WX4857,WX4786);
  not NOT_1591(WX4858,WX4857);
  not NOT_1592(WX4859,WX4787);
  not NOT_1593(WX4860,WX4859);
  not NOT_1594(WX4861,WX4788);
  not NOT_1595(WX4862,WX4861);
  not NOT_1596(WX4863,WX4789);
  not NOT_1597(WX4864,WX4863);
  not NOT_1598(WX4865,WX4790);
  not NOT_1599(WX4866,WX4865);
  not NOT_1600(WX4867,WX4791);
  not NOT_1601(WX4868,WX4867);
  not NOT_1602(WX4869,WX4792);
  not NOT_1603(WX4870,WX4869);
  not NOT_1604(WX4871,WX4793);
  not NOT_1605(WX4872,WX4871);
  not NOT_1606(WX4873,WX4794);
  not NOT_1607(WX4874,WX4873);
  not NOT_1608(WX4875,TM0);
  not NOT_1609(WX4876,TM0);
  not NOT_1610(WX4877,TM0);
  not NOT_1611(WX4878,TM1);
  not NOT_1612(WX4879,TM1);
  not NOT_1613(WX4880,WX4879);
  not NOT_1614(WX4881,WX4877);
  not NOT_1615(WX4882,WX4878);
  not NOT_1616(WX4883,WX4876);
  not NOT_1617(WX4884,WX4875);
  not NOT_1618(WX4888,WX4884);
  not NOT_1619(WX4890,WX4889);
  not NOT_1620(WX4891,WX4890);
  not NOT_1621(WX4895,WX4884);
  not NOT_1622(WX4897,WX4896);
  not NOT_1623(WX4898,WX4897);
  not NOT_1624(WX4902,WX4884);
  not NOT_1625(WX4904,WX4903);
  not NOT_1626(WX4905,WX4904);
  not NOT_1627(WX4909,WX4884);
  not NOT_1628(WX4911,WX4910);
  not NOT_1629(WX4912,WX4911);
  not NOT_1630(WX4916,WX4884);
  not NOT_1631(WX4918,WX4917);
  not NOT_1632(WX4919,WX4918);
  not NOT_1633(WX4923,WX4884);
  not NOT_1634(WX4925,WX4924);
  not NOT_1635(WX4926,WX4925);
  not NOT_1636(WX4930,WX4884);
  not NOT_1637(WX4932,WX4931);
  not NOT_1638(WX4933,WX4932);
  not NOT_1639(WX4937,WX4884);
  not NOT_1640(WX4939,WX4938);
  not NOT_1641(WX4940,WX4939);
  not NOT_1642(WX4944,WX4884);
  not NOT_1643(WX4946,WX4945);
  not NOT_1644(WX4947,WX4946);
  not NOT_1645(WX4951,WX4884);
  not NOT_1646(WX4953,WX4952);
  not NOT_1647(WX4954,WX4953);
  not NOT_1648(WX4958,WX4884);
  not NOT_1649(WX4960,WX4959);
  not NOT_1650(WX4961,WX4960);
  not NOT_1651(WX4965,WX4884);
  not NOT_1652(WX4967,WX4966);
  not NOT_1653(WX4968,WX4967);
  not NOT_1654(WX4972,WX4884);
  not NOT_1655(WX4974,WX4973);
  not NOT_1656(WX4975,WX4974);
  not NOT_1657(WX4979,WX4884);
  not NOT_1658(WX4981,WX4980);
  not NOT_1659(WX4982,WX4981);
  not NOT_1660(WX4986,WX4884);
  not NOT_1661(WX4988,WX4987);
  not NOT_1662(WX4989,WX4988);
  not NOT_1663(WX4993,WX4884);
  not NOT_1664(WX4995,WX4994);
  not NOT_1665(WX4996,WX4995);
  not NOT_1666(WX5000,WX4884);
  not NOT_1667(WX5002,WX5001);
  not NOT_1668(WX5003,WX5002);
  not NOT_1669(WX5007,WX4884);
  not NOT_1670(WX5009,WX5008);
  not NOT_1671(WX5010,WX5009);
  not NOT_1672(WX5014,WX4884);
  not NOT_1673(WX5016,WX5015);
  not NOT_1674(WX5017,WX5016);
  not NOT_1675(WX5021,WX4884);
  not NOT_1676(WX5023,WX5022);
  not NOT_1677(WX5024,WX5023);
  not NOT_1678(WX5028,WX4884);
  not NOT_1679(WX5030,WX5029);
  not NOT_1680(WX5031,WX5030);
  not NOT_1681(WX5035,WX4884);
  not NOT_1682(WX5037,WX5036);
  not NOT_1683(WX5038,WX5037);
  not NOT_1684(WX5042,WX4884);
  not NOT_1685(WX5044,WX5043);
  not NOT_1686(WX5045,WX5044);
  not NOT_1687(WX5049,WX4884);
  not NOT_1688(WX5051,WX5050);
  not NOT_1689(WX5052,WX5051);
  not NOT_1690(WX5056,WX4884);
  not NOT_1691(WX5058,WX5057);
  not NOT_1692(WX5059,WX5058);
  not NOT_1693(WX5063,WX4884);
  not NOT_1694(WX5065,WX5064);
  not NOT_1695(WX5066,WX5065);
  not NOT_1696(WX5070,WX4884);
  not NOT_1697(WX5072,WX5071);
  not NOT_1698(WX5073,WX5072);
  not NOT_1699(WX5077,WX4884);
  not NOT_1700(WX5079,WX5078);
  not NOT_1701(WX5080,WX5079);
  not NOT_1702(WX5084,WX4884);
  not NOT_1703(WX5086,WX5085);
  not NOT_1704(WX5087,WX5086);
  not NOT_1705(WX5091,WX4884);
  not NOT_1706(WX5093,WX5092);
  not NOT_1707(WX5094,WX5093);
  not NOT_1708(WX5098,WX4884);
  not NOT_1709(WX5100,WX5099);
  not NOT_1710(WX5101,WX5100);
  not NOT_1711(WX5105,WX4884);
  not NOT_1712(WX5107,WX5106);
  not NOT_1713(WX5108,WX5107);
  not NOT_1714(WX5109,RESET);
  not NOT_1715(WX5142,WX5109);
  not NOT_1716(WX5209,WX6175);
  not NOT_1717(WX5213,WX6176);
  not NOT_1718(WX5217,WX6176);
  not NOT_1719(WX5219,WX5210);
  not NOT_1720(WX5220,WX5219);
  not NOT_1721(WX5223,WX6175);
  not NOT_1722(WX5227,WX6176);
  not NOT_1723(WX5231,WX6176);
  not NOT_1724(WX5233,WX5224);
  not NOT_1725(WX5234,WX5233);
  not NOT_1726(WX5237,WX6175);
  not NOT_1727(WX5241,WX6176);
  not NOT_1728(WX5245,WX6176);
  not NOT_1729(WX5247,WX5238);
  not NOT_1730(WX5248,WX5247);
  not NOT_1731(WX5251,WX6175);
  not NOT_1732(WX5255,WX6176);
  not NOT_1733(WX5259,WX6176);
  not NOT_1734(WX5261,WX5252);
  not NOT_1735(WX5262,WX5261);
  not NOT_1736(WX5265,WX6175);
  not NOT_1737(WX5269,WX6176);
  not NOT_1738(WX5273,WX6176);
  not NOT_1739(WX5275,WX5266);
  not NOT_1740(WX5276,WX5275);
  not NOT_1741(WX5279,WX6175);
  not NOT_1742(WX5283,WX6176);
  not NOT_1743(WX5287,WX6176);
  not NOT_1744(WX5289,WX5280);
  not NOT_1745(WX5290,WX5289);
  not NOT_1746(WX5293,WX6175);
  not NOT_1747(WX5297,WX6176);
  not NOT_1748(WX5301,WX6176);
  not NOT_1749(WX5303,WX5294);
  not NOT_1750(WX5304,WX5303);
  not NOT_1751(WX5307,WX6175);
  not NOT_1752(WX5311,WX6176);
  not NOT_1753(WX5315,WX6176);
  not NOT_1754(WX5317,WX5308);
  not NOT_1755(WX5318,WX5317);
  not NOT_1756(WX5321,WX6175);
  not NOT_1757(WX5325,WX6176);
  not NOT_1758(WX5329,WX6176);
  not NOT_1759(WX5331,WX5322);
  not NOT_1760(WX5332,WX5331);
  not NOT_1761(WX5335,WX6175);
  not NOT_1762(WX5339,WX6176);
  not NOT_1763(WX5343,WX6176);
  not NOT_1764(WX5345,WX5336);
  not NOT_1765(WX5346,WX5345);
  not NOT_1766(WX5349,WX6175);
  not NOT_1767(WX5353,WX6176);
  not NOT_1768(WX5357,WX6176);
  not NOT_1769(WX5359,WX5350);
  not NOT_1770(WX5360,WX5359);
  not NOT_1771(WX5363,WX6175);
  not NOT_1772(WX5367,WX6176);
  not NOT_1773(WX5371,WX6176);
  not NOT_1774(WX5373,WX5364);
  not NOT_1775(WX5374,WX5373);
  not NOT_1776(WX5377,WX6175);
  not NOT_1777(WX5381,WX6176);
  not NOT_1778(WX5385,WX6176);
  not NOT_1779(WX5387,WX5378);
  not NOT_1780(WX5388,WX5387);
  not NOT_1781(WX5391,WX6175);
  not NOT_1782(WX5395,WX6176);
  not NOT_1783(WX5399,WX6176);
  not NOT_1784(WX5401,WX5392);
  not NOT_1785(WX5402,WX5401);
  not NOT_1786(WX5405,WX6175);
  not NOT_1787(WX5409,WX6176);
  not NOT_1788(WX5413,WX6176);
  not NOT_1789(WX5415,WX5406);
  not NOT_1790(WX5416,WX5415);
  not NOT_1791(WX5419,WX6175);
  not NOT_1792(WX5423,WX6176);
  not NOT_1793(WX5427,WX6176);
  not NOT_1794(WX5429,WX5420);
  not NOT_1795(WX5430,WX5429);
  not NOT_1796(WX5433,WX6175);
  not NOT_1797(WX5437,WX6176);
  not NOT_1798(WX5441,WX6176);
  not NOT_1799(WX5443,WX5434);
  not NOT_1800(WX5444,WX5443);
  not NOT_1801(WX5447,WX6175);
  not NOT_1802(WX5451,WX6176);
  not NOT_1803(WX5455,WX6176);
  not NOT_1804(WX5457,WX5448);
  not NOT_1805(WX5458,WX5457);
  not NOT_1806(WX5461,WX6175);
  not NOT_1807(WX5465,WX6176);
  not NOT_1808(WX5469,WX6176);
  not NOT_1809(WX5471,WX5462);
  not NOT_1810(WX5472,WX5471);
  not NOT_1811(WX5475,WX6175);
  not NOT_1812(WX5479,WX6176);
  not NOT_1813(WX5483,WX6176);
  not NOT_1814(WX5485,WX5476);
  not NOT_1815(WX5486,WX5485);
  not NOT_1816(WX5489,WX6175);
  not NOT_1817(WX5493,WX6176);
  not NOT_1818(WX5497,WX6176);
  not NOT_1819(WX5499,WX5490);
  not NOT_1820(WX5500,WX5499);
  not NOT_1821(WX5503,WX6175);
  not NOT_1822(WX5507,WX6176);
  not NOT_1823(WX5511,WX6176);
  not NOT_1824(WX5513,WX5504);
  not NOT_1825(WX5514,WX5513);
  not NOT_1826(WX5517,WX6175);
  not NOT_1827(WX5521,WX6176);
  not NOT_1828(WX5525,WX6176);
  not NOT_1829(WX5527,WX5518);
  not NOT_1830(WX5528,WX5527);
  not NOT_1831(WX5531,WX6175);
  not NOT_1832(WX5535,WX6176);
  not NOT_1833(WX5539,WX6176);
  not NOT_1834(WX5541,WX5532);
  not NOT_1835(WX5542,WX5541);
  not NOT_1836(WX5545,WX6175);
  not NOT_1837(WX5549,WX6176);
  not NOT_1838(WX5553,WX6176);
  not NOT_1839(WX5555,WX5546);
  not NOT_1840(WX5556,WX5555);
  not NOT_1841(WX5559,WX6175);
  not NOT_1842(WX5563,WX6176);
  not NOT_1843(WX5567,WX6176);
  not NOT_1844(WX5569,WX5560);
  not NOT_1845(WX5570,WX5569);
  not NOT_1846(WX5573,WX6175);
  not NOT_1847(WX5577,WX6176);
  not NOT_1848(WX5581,WX6176);
  not NOT_1849(WX5583,WX5574);
  not NOT_1850(WX5584,WX5583);
  not NOT_1851(WX5587,WX6175);
  not NOT_1852(WX5591,WX6176);
  not NOT_1853(WX5595,WX6176);
  not NOT_1854(WX5597,WX5588);
  not NOT_1855(WX5598,WX5597);
  not NOT_1856(WX5601,WX6175);
  not NOT_1857(WX5605,WX6176);
  not NOT_1858(WX5609,WX6176);
  not NOT_1859(WX5611,WX5602);
  not NOT_1860(WX5612,WX5611);
  not NOT_1861(WX5615,WX6175);
  not NOT_1862(WX5619,WX6176);
  not NOT_1863(WX5623,WX6176);
  not NOT_1864(WX5625,WX5616);
  not NOT_1865(WX5626,WX5625);
  not NOT_1866(WX5629,WX6175);
  not NOT_1867(WX5633,WX6176);
  not NOT_1868(WX5637,WX6176);
  not NOT_1869(WX5639,WX5630);
  not NOT_1870(WX5640,WX5639);
  not NOT_1871(WX5643,WX6175);
  not NOT_1872(WX5647,WX6176);
  not NOT_1873(WX5651,WX6176);
  not NOT_1874(WX5653,WX5644);
  not NOT_1875(WX5654,WX5653);
  not NOT_1876(WX5655,WX5657);
  not NOT_1877(WX5720,WX6137);
  not NOT_1878(WX5721,WX6139);
  not NOT_1879(WX5722,WX6141);
  not NOT_1880(WX5723,WX6143);
  not NOT_1881(WX5724,WX6145);
  not NOT_1882(WX5725,WX6147);
  not NOT_1883(WX5726,WX6149);
  not NOT_1884(WX5727,WX6151);
  not NOT_1885(WX5728,WX6153);
  not NOT_1886(WX5729,WX6155);
  not NOT_1887(WX5730,WX6157);
  not NOT_1888(WX5731,WX6159);
  not NOT_1889(WX5732,WX6161);
  not NOT_1890(WX5733,WX6163);
  not NOT_1891(WX5734,WX6165);
  not NOT_1892(WX5735,WX6167);
  not NOT_1893(WX5736,WX6105);
  not NOT_1894(WX5737,WX6107);
  not NOT_1895(WX5738,WX6109);
  not NOT_1896(WX5739,WX6111);
  not NOT_1897(WX5740,WX6113);
  not NOT_1898(WX5741,WX6115);
  not NOT_1899(WX5742,WX6117);
  not NOT_1900(WX5743,WX6119);
  not NOT_1901(WX5744,WX6121);
  not NOT_1902(WX5745,WX6123);
  not NOT_1903(WX5746,WX6125);
  not NOT_1904(WX5747,WX6127);
  not NOT_1905(WX5748,WX6129);
  not NOT_1906(WX5749,WX6131);
  not NOT_1907(WX5750,WX6133);
  not NOT_1908(WX5751,WX6135);
  not NOT_1909(WX5752,WX5720);
  not NOT_1910(WX5753,WX5721);
  not NOT_1911(WX5754,WX5722);
  not NOT_1912(WX5755,WX5723);
  not NOT_1913(WX5756,WX5724);
  not NOT_1914(WX5757,WX5725);
  not NOT_1915(WX5758,WX5726);
  not NOT_1916(WX5759,WX5727);
  not NOT_1917(WX5760,WX5728);
  not NOT_1918(WX5761,WX5729);
  not NOT_1919(WX5762,WX5730);
  not NOT_1920(WX5763,WX5731);
  not NOT_1921(WX5764,WX5732);
  not NOT_1922(WX5765,WX5733);
  not NOT_1923(WX5766,WX5734);
  not NOT_1924(WX5767,WX5735);
  not NOT_1925(WX5768,WX5736);
  not NOT_1926(WX5769,WX5737);
  not NOT_1927(WX5770,WX5738);
  not NOT_1928(WX5771,WX5739);
  not NOT_1929(WX5772,WX5740);
  not NOT_1930(WX5773,WX5741);
  not NOT_1931(WX5774,WX5742);
  not NOT_1932(WX5775,WX5743);
  not NOT_1933(WX5776,WX5744);
  not NOT_1934(WX5777,WX5745);
  not NOT_1935(WX5778,WX5746);
  not NOT_1936(WX5779,WX5747);
  not NOT_1937(WX5780,WX5748);
  not NOT_1938(WX5781,WX5749);
  not NOT_1939(WX5782,WX5750);
  not NOT_1940(WX5783,WX5751);
  not NOT_1941(WX5784,WX6009);
  not NOT_1942(WX5785,WX6011);
  not NOT_1943(WX5786,WX6013);
  not NOT_1944(WX5787,WX6015);
  not NOT_1945(WX5788,WX6017);
  not NOT_1946(WX5789,WX6019);
  not NOT_1947(WX5790,WX6021);
  not NOT_1948(WX5791,WX6023);
  not NOT_1949(WX5792,WX6025);
  not NOT_1950(WX5793,WX6027);
  not NOT_1951(WX5794,WX6029);
  not NOT_1952(WX5795,WX6031);
  not NOT_1953(WX5796,WX6033);
  not NOT_1954(WX5797,WX6035);
  not NOT_1955(WX5798,WX6037);
  not NOT_1956(WX5799,WX6039);
  not NOT_1957(WX5800,WX6041);
  not NOT_1958(WX5801,WX6043);
  not NOT_1959(WX5802,WX6045);
  not NOT_1960(WX5803,WX6047);
  not NOT_1961(WX5804,WX6049);
  not NOT_1962(WX5805,WX6051);
  not NOT_1963(WX5806,WX6053);
  not NOT_1964(WX5807,WX6055);
  not NOT_1965(WX5808,WX6057);
  not NOT_1966(WX5809,WX6059);
  not NOT_1967(WX5810,WX6061);
  not NOT_1968(WX5811,WX6063);
  not NOT_1969(WX5812,WX6065);
  not NOT_1970(WX5813,WX6067);
  not NOT_1971(WX5814,WX6069);
  not NOT_1972(WX5815,WX6071);
  not NOT_1973(WX6104,WX6088);
  not NOT_1974(WX6105,WX6104);
  not NOT_1975(WX6106,WX6089);
  not NOT_1976(WX6107,WX6106);
  not NOT_1977(WX6108,WX6090);
  not NOT_1978(WX6109,WX6108);
  not NOT_1979(WX6110,WX6091);
  not NOT_1980(WX6111,WX6110);
  not NOT_1981(WX6112,WX6092);
  not NOT_1982(WX6113,WX6112);
  not NOT_1983(WX6114,WX6093);
  not NOT_1984(WX6115,WX6114);
  not NOT_1985(WX6116,WX6094);
  not NOT_1986(WX6117,WX6116);
  not NOT_1987(WX6118,WX6095);
  not NOT_1988(WX6119,WX6118);
  not NOT_1989(WX6120,WX6096);
  not NOT_1990(WX6121,WX6120);
  not NOT_1991(WX6122,WX6097);
  not NOT_1992(WX6123,WX6122);
  not NOT_1993(WX6124,WX6098);
  not NOT_1994(WX6125,WX6124);
  not NOT_1995(WX6126,WX6099);
  not NOT_1996(WX6127,WX6126);
  not NOT_1997(WX6128,WX6100);
  not NOT_1998(WX6129,WX6128);
  not NOT_1999(WX6130,WX6101);
  not NOT_2000(WX6131,WX6130);
  not NOT_2001(WX6132,WX6102);
  not NOT_2002(WX6133,WX6132);
  not NOT_2003(WX6134,WX6103);
  not NOT_2004(WX6135,WX6134);
  not NOT_2005(WX6136,WX6072);
  not NOT_2006(WX6137,WX6136);
  not NOT_2007(WX6138,WX6073);
  not NOT_2008(WX6139,WX6138);
  not NOT_2009(WX6140,WX6074);
  not NOT_2010(WX6141,WX6140);
  not NOT_2011(WX6142,WX6075);
  not NOT_2012(WX6143,WX6142);
  not NOT_2013(WX6144,WX6076);
  not NOT_2014(WX6145,WX6144);
  not NOT_2015(WX6146,WX6077);
  not NOT_2016(WX6147,WX6146);
  not NOT_2017(WX6148,WX6078);
  not NOT_2018(WX6149,WX6148);
  not NOT_2019(WX6150,WX6079);
  not NOT_2020(WX6151,WX6150);
  not NOT_2021(WX6152,WX6080);
  not NOT_2022(WX6153,WX6152);
  not NOT_2023(WX6154,WX6081);
  not NOT_2024(WX6155,WX6154);
  not NOT_2025(WX6156,WX6082);
  not NOT_2026(WX6157,WX6156);
  not NOT_2027(WX6158,WX6083);
  not NOT_2028(WX6159,WX6158);
  not NOT_2029(WX6160,WX6084);
  not NOT_2030(WX6161,WX6160);
  not NOT_2031(WX6162,WX6085);
  not NOT_2032(WX6163,WX6162);
  not NOT_2033(WX6164,WX6086);
  not NOT_2034(WX6165,WX6164);
  not NOT_2035(WX6166,WX6087);
  not NOT_2036(WX6167,WX6166);
  not NOT_2037(WX6168,TM0);
  not NOT_2038(WX6169,TM0);
  not NOT_2039(WX6170,TM0);
  not NOT_2040(WX6171,TM1);
  not NOT_2041(WX6172,TM1);
  not NOT_2042(WX6173,WX6172);
  not NOT_2043(WX6174,WX6170);
  not NOT_2044(WX6175,WX6171);
  not NOT_2045(WX6176,WX6169);
  not NOT_2046(WX6177,WX6168);
  not NOT_2047(WX6181,WX6177);
  not NOT_2048(WX6183,WX6182);
  not NOT_2049(WX6184,WX6183);
  not NOT_2050(WX6188,WX6177);
  not NOT_2051(WX6190,WX6189);
  not NOT_2052(WX6191,WX6190);
  not NOT_2053(WX6195,WX6177);
  not NOT_2054(WX6197,WX6196);
  not NOT_2055(WX6198,WX6197);
  not NOT_2056(WX6202,WX6177);
  not NOT_2057(WX6204,WX6203);
  not NOT_2058(WX6205,WX6204);
  not NOT_2059(WX6209,WX6177);
  not NOT_2060(WX6211,WX6210);
  not NOT_2061(WX6212,WX6211);
  not NOT_2062(WX6216,WX6177);
  not NOT_2063(WX6218,WX6217);
  not NOT_2064(WX6219,WX6218);
  not NOT_2065(WX6223,WX6177);
  not NOT_2066(WX6225,WX6224);
  not NOT_2067(WX6226,WX6225);
  not NOT_2068(WX6230,WX6177);
  not NOT_2069(WX6232,WX6231);
  not NOT_2070(WX6233,WX6232);
  not NOT_2071(WX6237,WX6177);
  not NOT_2072(WX6239,WX6238);
  not NOT_2073(WX6240,WX6239);
  not NOT_2074(WX6244,WX6177);
  not NOT_2075(WX6246,WX6245);
  not NOT_2076(WX6247,WX6246);
  not NOT_2077(WX6251,WX6177);
  not NOT_2078(WX6253,WX6252);
  not NOT_2079(WX6254,WX6253);
  not NOT_2080(WX6258,WX6177);
  not NOT_2081(WX6260,WX6259);
  not NOT_2082(WX6261,WX6260);
  not NOT_2083(WX6265,WX6177);
  not NOT_2084(WX6267,WX6266);
  not NOT_2085(WX6268,WX6267);
  not NOT_2086(WX6272,WX6177);
  not NOT_2087(WX6274,WX6273);
  not NOT_2088(WX6275,WX6274);
  not NOT_2089(WX6279,WX6177);
  not NOT_2090(WX6281,WX6280);
  not NOT_2091(WX6282,WX6281);
  not NOT_2092(WX6286,WX6177);
  not NOT_2093(WX6288,WX6287);
  not NOT_2094(WX6289,WX6288);
  not NOT_2095(WX6293,WX6177);
  not NOT_2096(WX6295,WX6294);
  not NOT_2097(WX6296,WX6295);
  not NOT_2098(WX6300,WX6177);
  not NOT_2099(WX6302,WX6301);
  not NOT_2100(WX6303,WX6302);
  not NOT_2101(WX6307,WX6177);
  not NOT_2102(WX6309,WX6308);
  not NOT_2103(WX6310,WX6309);
  not NOT_2104(WX6314,WX6177);
  not NOT_2105(WX6316,WX6315);
  not NOT_2106(WX6317,WX6316);
  not NOT_2107(WX6321,WX6177);
  not NOT_2108(WX6323,WX6322);
  not NOT_2109(WX6324,WX6323);
  not NOT_2110(WX6328,WX6177);
  not NOT_2111(WX6330,WX6329);
  not NOT_2112(WX6331,WX6330);
  not NOT_2113(WX6335,WX6177);
  not NOT_2114(WX6337,WX6336);
  not NOT_2115(WX6338,WX6337);
  not NOT_2116(WX6342,WX6177);
  not NOT_2117(WX6344,WX6343);
  not NOT_2118(WX6345,WX6344);
  not NOT_2119(WX6349,WX6177);
  not NOT_2120(WX6351,WX6350);
  not NOT_2121(WX6352,WX6351);
  not NOT_2122(WX6356,WX6177);
  not NOT_2123(WX6358,WX6357);
  not NOT_2124(WX6359,WX6358);
  not NOT_2125(WX6363,WX6177);
  not NOT_2126(WX6365,WX6364);
  not NOT_2127(WX6366,WX6365);
  not NOT_2128(WX6370,WX6177);
  not NOT_2129(WX6372,WX6371);
  not NOT_2130(WX6373,WX6372);
  not NOT_2131(WX6377,WX6177);
  not NOT_2132(WX6379,WX6378);
  not NOT_2133(WX6380,WX6379);
  not NOT_2134(WX6384,WX6177);
  not NOT_2135(WX6386,WX6385);
  not NOT_2136(WX6387,WX6386);
  not NOT_2137(WX6391,WX6177);
  not NOT_2138(WX6393,WX6392);
  not NOT_2139(WX6394,WX6393);
  not NOT_2140(WX6398,WX6177);
  not NOT_2141(WX6400,WX6399);
  not NOT_2142(WX6401,WX6400);
  not NOT_2143(WX6402,RESET);
  not NOT_2144(WX6435,WX6402);
  not NOT_2145(WX6502,WX7468);
  not NOT_2146(WX6506,WX7469);
  not NOT_2147(WX6510,WX7469);
  not NOT_2148(WX6512,WX6503);
  not NOT_2149(WX6513,WX6512);
  not NOT_2150(WX6516,WX7468);
  not NOT_2151(WX6520,WX7469);
  not NOT_2152(WX6524,WX7469);
  not NOT_2153(WX6526,WX6517);
  not NOT_2154(WX6527,WX6526);
  not NOT_2155(WX6530,WX7468);
  not NOT_2156(WX6534,WX7469);
  not NOT_2157(WX6538,WX7469);
  not NOT_2158(WX6540,WX6531);
  not NOT_2159(WX6541,WX6540);
  not NOT_2160(WX6544,WX7468);
  not NOT_2161(WX6548,WX7469);
  not NOT_2162(WX6552,WX7469);
  not NOT_2163(WX6554,WX6545);
  not NOT_2164(WX6555,WX6554);
  not NOT_2165(WX6558,WX7468);
  not NOT_2166(WX6562,WX7469);
  not NOT_2167(WX6566,WX7469);
  not NOT_2168(WX6568,WX6559);
  not NOT_2169(WX6569,WX6568);
  not NOT_2170(WX6572,WX7468);
  not NOT_2171(WX6576,WX7469);
  not NOT_2172(WX6580,WX7469);
  not NOT_2173(WX6582,WX6573);
  not NOT_2174(WX6583,WX6582);
  not NOT_2175(WX6586,WX7468);
  not NOT_2176(WX6590,WX7469);
  not NOT_2177(WX6594,WX7469);
  not NOT_2178(WX6596,WX6587);
  not NOT_2179(WX6597,WX6596);
  not NOT_2180(WX6600,WX7468);
  not NOT_2181(WX6604,WX7469);
  not NOT_2182(WX6608,WX7469);
  not NOT_2183(WX6610,WX6601);
  not NOT_2184(WX6611,WX6610);
  not NOT_2185(WX6614,WX7468);
  not NOT_2186(WX6618,WX7469);
  not NOT_2187(WX6622,WX7469);
  not NOT_2188(WX6624,WX6615);
  not NOT_2189(WX6625,WX6624);
  not NOT_2190(WX6628,WX7468);
  not NOT_2191(WX6632,WX7469);
  not NOT_2192(WX6636,WX7469);
  not NOT_2193(WX6638,WX6629);
  not NOT_2194(WX6639,WX6638);
  not NOT_2195(WX6642,WX7468);
  not NOT_2196(WX6646,WX7469);
  not NOT_2197(WX6650,WX7469);
  not NOT_2198(WX6652,WX6643);
  not NOT_2199(WX6653,WX6652);
  not NOT_2200(WX6656,WX7468);
  not NOT_2201(WX6660,WX7469);
  not NOT_2202(WX6664,WX7469);
  not NOT_2203(WX6666,WX6657);
  not NOT_2204(WX6667,WX6666);
  not NOT_2205(WX6670,WX7468);
  not NOT_2206(WX6674,WX7469);
  not NOT_2207(WX6678,WX7469);
  not NOT_2208(WX6680,WX6671);
  not NOT_2209(WX6681,WX6680);
  not NOT_2210(WX6684,WX7468);
  not NOT_2211(WX6688,WX7469);
  not NOT_2212(WX6692,WX7469);
  not NOT_2213(WX6694,WX6685);
  not NOT_2214(WX6695,WX6694);
  not NOT_2215(WX6698,WX7468);
  not NOT_2216(WX6702,WX7469);
  not NOT_2217(WX6706,WX7469);
  not NOT_2218(WX6708,WX6699);
  not NOT_2219(WX6709,WX6708);
  not NOT_2220(WX6712,WX7468);
  not NOT_2221(WX6716,WX7469);
  not NOT_2222(WX6720,WX7469);
  not NOT_2223(WX6722,WX6713);
  not NOT_2224(WX6723,WX6722);
  not NOT_2225(WX6726,WX7468);
  not NOT_2226(WX6730,WX7469);
  not NOT_2227(WX6734,WX7469);
  not NOT_2228(WX6736,WX6727);
  not NOT_2229(WX6737,WX6736);
  not NOT_2230(WX6740,WX7468);
  not NOT_2231(WX6744,WX7469);
  not NOT_2232(WX6748,WX7469);
  not NOT_2233(WX6750,WX6741);
  not NOT_2234(WX6751,WX6750);
  not NOT_2235(WX6754,WX7468);
  not NOT_2236(WX6758,WX7469);
  not NOT_2237(WX6762,WX7469);
  not NOT_2238(WX6764,WX6755);
  not NOT_2239(WX6765,WX6764);
  not NOT_2240(WX6768,WX7468);
  not NOT_2241(WX6772,WX7469);
  not NOT_2242(WX6776,WX7469);
  not NOT_2243(WX6778,WX6769);
  not NOT_2244(WX6779,WX6778);
  not NOT_2245(WX6782,WX7468);
  not NOT_2246(WX6786,WX7469);
  not NOT_2247(WX6790,WX7469);
  not NOT_2248(WX6792,WX6783);
  not NOT_2249(WX6793,WX6792);
  not NOT_2250(WX6796,WX7468);
  not NOT_2251(WX6800,WX7469);
  not NOT_2252(WX6804,WX7469);
  not NOT_2253(WX6806,WX6797);
  not NOT_2254(WX6807,WX6806);
  not NOT_2255(WX6810,WX7468);
  not NOT_2256(WX6814,WX7469);
  not NOT_2257(WX6818,WX7469);
  not NOT_2258(WX6820,WX6811);
  not NOT_2259(WX6821,WX6820);
  not NOT_2260(WX6824,WX7468);
  not NOT_2261(WX6828,WX7469);
  not NOT_2262(WX6832,WX7469);
  not NOT_2263(WX6834,WX6825);
  not NOT_2264(WX6835,WX6834);
  not NOT_2265(WX6838,WX7468);
  not NOT_2266(WX6842,WX7469);
  not NOT_2267(WX6846,WX7469);
  not NOT_2268(WX6848,WX6839);
  not NOT_2269(WX6849,WX6848);
  not NOT_2270(WX6852,WX7468);
  not NOT_2271(WX6856,WX7469);
  not NOT_2272(WX6860,WX7469);
  not NOT_2273(WX6862,WX6853);
  not NOT_2274(WX6863,WX6862);
  not NOT_2275(WX6866,WX7468);
  not NOT_2276(WX6870,WX7469);
  not NOT_2277(WX6874,WX7469);
  not NOT_2278(WX6876,WX6867);
  not NOT_2279(WX6877,WX6876);
  not NOT_2280(WX6880,WX7468);
  not NOT_2281(WX6884,WX7469);
  not NOT_2282(WX6888,WX7469);
  not NOT_2283(WX6890,WX6881);
  not NOT_2284(WX6891,WX6890);
  not NOT_2285(WX6894,WX7468);
  not NOT_2286(WX6898,WX7469);
  not NOT_2287(WX6902,WX7469);
  not NOT_2288(WX6904,WX6895);
  not NOT_2289(WX6905,WX6904);
  not NOT_2290(WX6908,WX7468);
  not NOT_2291(WX6912,WX7469);
  not NOT_2292(WX6916,WX7469);
  not NOT_2293(WX6918,WX6909);
  not NOT_2294(WX6919,WX6918);
  not NOT_2295(WX6922,WX7468);
  not NOT_2296(WX6926,WX7469);
  not NOT_2297(WX6930,WX7469);
  not NOT_2298(WX6932,WX6923);
  not NOT_2299(WX6933,WX6932);
  not NOT_2300(WX6936,WX7468);
  not NOT_2301(WX6940,WX7469);
  not NOT_2302(WX6944,WX7469);
  not NOT_2303(WX6946,WX6937);
  not NOT_2304(WX6947,WX6946);
  not NOT_2305(WX6948,WX6950);
  not NOT_2306(WX7013,WX7430);
  not NOT_2307(WX7014,WX7432);
  not NOT_2308(WX7015,WX7434);
  not NOT_2309(WX7016,WX7436);
  not NOT_2310(WX7017,WX7438);
  not NOT_2311(WX7018,WX7440);
  not NOT_2312(WX7019,WX7442);
  not NOT_2313(WX7020,WX7444);
  not NOT_2314(WX7021,WX7446);
  not NOT_2315(WX7022,WX7448);
  not NOT_2316(WX7023,WX7450);
  not NOT_2317(WX7024,WX7452);
  not NOT_2318(WX7025,WX7454);
  not NOT_2319(WX7026,WX7456);
  not NOT_2320(WX7027,WX7458);
  not NOT_2321(WX7028,WX7460);
  not NOT_2322(WX7029,WX7398);
  not NOT_2323(WX7030,WX7400);
  not NOT_2324(WX7031,WX7402);
  not NOT_2325(WX7032,WX7404);
  not NOT_2326(WX7033,WX7406);
  not NOT_2327(WX7034,WX7408);
  not NOT_2328(WX7035,WX7410);
  not NOT_2329(WX7036,WX7412);
  not NOT_2330(WX7037,WX7414);
  not NOT_2331(WX7038,WX7416);
  not NOT_2332(WX7039,WX7418);
  not NOT_2333(WX7040,WX7420);
  not NOT_2334(WX7041,WX7422);
  not NOT_2335(WX7042,WX7424);
  not NOT_2336(WX7043,WX7426);
  not NOT_2337(WX7044,WX7428);
  not NOT_2338(WX7045,WX7013);
  not NOT_2339(WX7046,WX7014);
  not NOT_2340(WX7047,WX7015);
  not NOT_2341(WX7048,WX7016);
  not NOT_2342(WX7049,WX7017);
  not NOT_2343(WX7050,WX7018);
  not NOT_2344(WX7051,WX7019);
  not NOT_2345(WX7052,WX7020);
  not NOT_2346(WX7053,WX7021);
  not NOT_2347(WX7054,WX7022);
  not NOT_2348(WX7055,WX7023);
  not NOT_2349(WX7056,WX7024);
  not NOT_2350(WX7057,WX7025);
  not NOT_2351(WX7058,WX7026);
  not NOT_2352(WX7059,WX7027);
  not NOT_2353(WX7060,WX7028);
  not NOT_2354(WX7061,WX7029);
  not NOT_2355(WX7062,WX7030);
  not NOT_2356(WX7063,WX7031);
  not NOT_2357(WX7064,WX7032);
  not NOT_2358(WX7065,WX7033);
  not NOT_2359(WX7066,WX7034);
  not NOT_2360(WX7067,WX7035);
  not NOT_2361(WX7068,WX7036);
  not NOT_2362(WX7069,WX7037);
  not NOT_2363(WX7070,WX7038);
  not NOT_2364(WX7071,WX7039);
  not NOT_2365(WX7072,WX7040);
  not NOT_2366(WX7073,WX7041);
  not NOT_2367(WX7074,WX7042);
  not NOT_2368(WX7075,WX7043);
  not NOT_2369(WX7076,WX7044);
  not NOT_2370(WX7077,WX7302);
  not NOT_2371(WX7078,WX7304);
  not NOT_2372(WX7079,WX7306);
  not NOT_2373(WX7080,WX7308);
  not NOT_2374(WX7081,WX7310);
  not NOT_2375(WX7082,WX7312);
  not NOT_2376(WX7083,WX7314);
  not NOT_2377(WX7084,WX7316);
  not NOT_2378(WX7085,WX7318);
  not NOT_2379(WX7086,WX7320);
  not NOT_2380(WX7087,WX7322);
  not NOT_2381(WX7088,WX7324);
  not NOT_2382(WX7089,WX7326);
  not NOT_2383(WX7090,WX7328);
  not NOT_2384(WX7091,WX7330);
  not NOT_2385(WX7092,WX7332);
  not NOT_2386(WX7093,WX7334);
  not NOT_2387(WX7094,WX7336);
  not NOT_2388(WX7095,WX7338);
  not NOT_2389(WX7096,WX7340);
  not NOT_2390(WX7097,WX7342);
  not NOT_2391(WX7098,WX7344);
  not NOT_2392(WX7099,WX7346);
  not NOT_2393(WX7100,WX7348);
  not NOT_2394(WX7101,WX7350);
  not NOT_2395(WX7102,WX7352);
  not NOT_2396(WX7103,WX7354);
  not NOT_2397(WX7104,WX7356);
  not NOT_2398(WX7105,WX7358);
  not NOT_2399(WX7106,WX7360);
  not NOT_2400(WX7107,WX7362);
  not NOT_2401(WX7108,WX7364);
  not NOT_2402(WX7397,WX7381);
  not NOT_2403(WX7398,WX7397);
  not NOT_2404(WX7399,WX7382);
  not NOT_2405(WX7400,WX7399);
  not NOT_2406(WX7401,WX7383);
  not NOT_2407(WX7402,WX7401);
  not NOT_2408(WX7403,WX7384);
  not NOT_2409(WX7404,WX7403);
  not NOT_2410(WX7405,WX7385);
  not NOT_2411(WX7406,WX7405);
  not NOT_2412(WX7407,WX7386);
  not NOT_2413(WX7408,WX7407);
  not NOT_2414(WX7409,WX7387);
  not NOT_2415(WX7410,WX7409);
  not NOT_2416(WX7411,WX7388);
  not NOT_2417(WX7412,WX7411);
  not NOT_2418(WX7413,WX7389);
  not NOT_2419(WX7414,WX7413);
  not NOT_2420(WX7415,WX7390);
  not NOT_2421(WX7416,WX7415);
  not NOT_2422(WX7417,WX7391);
  not NOT_2423(WX7418,WX7417);
  not NOT_2424(WX7419,WX7392);
  not NOT_2425(WX7420,WX7419);
  not NOT_2426(WX7421,WX7393);
  not NOT_2427(WX7422,WX7421);
  not NOT_2428(WX7423,WX7394);
  not NOT_2429(WX7424,WX7423);
  not NOT_2430(WX7425,WX7395);
  not NOT_2431(WX7426,WX7425);
  not NOT_2432(WX7427,WX7396);
  not NOT_2433(WX7428,WX7427);
  not NOT_2434(WX7429,WX7365);
  not NOT_2435(WX7430,WX7429);
  not NOT_2436(WX7431,WX7366);
  not NOT_2437(WX7432,WX7431);
  not NOT_2438(WX7433,WX7367);
  not NOT_2439(WX7434,WX7433);
  not NOT_2440(WX7435,WX7368);
  not NOT_2441(WX7436,WX7435);
  not NOT_2442(WX7437,WX7369);
  not NOT_2443(WX7438,WX7437);
  not NOT_2444(WX7439,WX7370);
  not NOT_2445(WX7440,WX7439);
  not NOT_2446(WX7441,WX7371);
  not NOT_2447(WX7442,WX7441);
  not NOT_2448(WX7443,WX7372);
  not NOT_2449(WX7444,WX7443);
  not NOT_2450(WX7445,WX7373);
  not NOT_2451(WX7446,WX7445);
  not NOT_2452(WX7447,WX7374);
  not NOT_2453(WX7448,WX7447);
  not NOT_2454(WX7449,WX7375);
  not NOT_2455(WX7450,WX7449);
  not NOT_2456(WX7451,WX7376);
  not NOT_2457(WX7452,WX7451);
  not NOT_2458(WX7453,WX7377);
  not NOT_2459(WX7454,WX7453);
  not NOT_2460(WX7455,WX7378);
  not NOT_2461(WX7456,WX7455);
  not NOT_2462(WX7457,WX7379);
  not NOT_2463(WX7458,WX7457);
  not NOT_2464(WX7459,WX7380);
  not NOT_2465(WX7460,WX7459);
  not NOT_2466(WX7461,TM0);
  not NOT_2467(WX7462,TM0);
  not NOT_2468(WX7463,TM0);
  not NOT_2469(WX7464,TM1);
  not NOT_2470(WX7465,TM1);
  not NOT_2471(WX7466,WX7465);
  not NOT_2472(WX7467,WX7463);
  not NOT_2473(WX7468,WX7464);
  not NOT_2474(WX7469,WX7462);
  not NOT_2475(WX7470,WX7461);
  not NOT_2476(WX7474,WX7470);
  not NOT_2477(WX7476,WX7475);
  not NOT_2478(WX7477,WX7476);
  not NOT_2479(WX7481,WX7470);
  not NOT_2480(WX7483,WX7482);
  not NOT_2481(WX7484,WX7483);
  not NOT_2482(WX7488,WX7470);
  not NOT_2483(WX7490,WX7489);
  not NOT_2484(WX7491,WX7490);
  not NOT_2485(WX7495,WX7470);
  not NOT_2486(WX7497,WX7496);
  not NOT_2487(WX7498,WX7497);
  not NOT_2488(WX7502,WX7470);
  not NOT_2489(WX7504,WX7503);
  not NOT_2490(WX7505,WX7504);
  not NOT_2491(WX7509,WX7470);
  not NOT_2492(WX7511,WX7510);
  not NOT_2493(WX7512,WX7511);
  not NOT_2494(WX7516,WX7470);
  not NOT_2495(WX7518,WX7517);
  not NOT_2496(WX7519,WX7518);
  not NOT_2497(WX7523,WX7470);
  not NOT_2498(WX7525,WX7524);
  not NOT_2499(WX7526,WX7525);
  not NOT_2500(WX7530,WX7470);
  not NOT_2501(WX7532,WX7531);
  not NOT_2502(WX7533,WX7532);
  not NOT_2503(WX7537,WX7470);
  not NOT_2504(WX7539,WX7538);
  not NOT_2505(WX7540,WX7539);
  not NOT_2506(WX7544,WX7470);
  not NOT_2507(WX7546,WX7545);
  not NOT_2508(WX7547,WX7546);
  not NOT_2509(WX7551,WX7470);
  not NOT_2510(WX7553,WX7552);
  not NOT_2511(WX7554,WX7553);
  not NOT_2512(WX7558,WX7470);
  not NOT_2513(WX7560,WX7559);
  not NOT_2514(WX7561,WX7560);
  not NOT_2515(WX7565,WX7470);
  not NOT_2516(WX7567,WX7566);
  not NOT_2517(WX7568,WX7567);
  not NOT_2518(WX7572,WX7470);
  not NOT_2519(WX7574,WX7573);
  not NOT_2520(WX7575,WX7574);
  not NOT_2521(WX7579,WX7470);
  not NOT_2522(WX7581,WX7580);
  not NOT_2523(WX7582,WX7581);
  not NOT_2524(WX7586,WX7470);
  not NOT_2525(WX7588,WX7587);
  not NOT_2526(WX7589,WX7588);
  not NOT_2527(WX7593,WX7470);
  not NOT_2528(WX7595,WX7594);
  not NOT_2529(WX7596,WX7595);
  not NOT_2530(WX7600,WX7470);
  not NOT_2531(WX7602,WX7601);
  not NOT_2532(WX7603,WX7602);
  not NOT_2533(WX7607,WX7470);
  not NOT_2534(WX7609,WX7608);
  not NOT_2535(WX7610,WX7609);
  not NOT_2536(WX7614,WX7470);
  not NOT_2537(WX7616,WX7615);
  not NOT_2538(WX7617,WX7616);
  not NOT_2539(WX7621,WX7470);
  not NOT_2540(WX7623,WX7622);
  not NOT_2541(WX7624,WX7623);
  not NOT_2542(WX7628,WX7470);
  not NOT_2543(WX7630,WX7629);
  not NOT_2544(WX7631,WX7630);
  not NOT_2545(WX7635,WX7470);
  not NOT_2546(WX7637,WX7636);
  not NOT_2547(WX7638,WX7637);
  not NOT_2548(WX7642,WX7470);
  not NOT_2549(WX7644,WX7643);
  not NOT_2550(WX7645,WX7644);
  not NOT_2551(WX7649,WX7470);
  not NOT_2552(WX7651,WX7650);
  not NOT_2553(WX7652,WX7651);
  not NOT_2554(WX7656,WX7470);
  not NOT_2555(WX7658,WX7657);
  not NOT_2556(WX7659,WX7658);
  not NOT_2557(WX7663,WX7470);
  not NOT_2558(WX7665,WX7664);
  not NOT_2559(WX7666,WX7665);
  not NOT_2560(WX7670,WX7470);
  not NOT_2561(WX7672,WX7671);
  not NOT_2562(WX7673,WX7672);
  not NOT_2563(WX7677,WX7470);
  not NOT_2564(WX7679,WX7678);
  not NOT_2565(WX7680,WX7679);
  not NOT_2566(WX7684,WX7470);
  not NOT_2567(WX7686,WX7685);
  not NOT_2568(WX7687,WX7686);
  not NOT_2569(WX7691,WX7470);
  not NOT_2570(WX7693,WX7692);
  not NOT_2571(WX7694,WX7693);
  not NOT_2572(WX7695,RESET);
  not NOT_2573(WX7728,WX7695);
  not NOT_2574(WX7795,WX8761);
  not NOT_2575(WX7799,WX8762);
  not NOT_2576(WX7803,WX8762);
  not NOT_2577(WX7805,WX7796);
  not NOT_2578(WX7806,WX7805);
  not NOT_2579(WX7809,WX8761);
  not NOT_2580(WX7813,WX8762);
  not NOT_2581(WX7817,WX8762);
  not NOT_2582(WX7819,WX7810);
  not NOT_2583(WX7820,WX7819);
  not NOT_2584(WX7823,WX8761);
  not NOT_2585(WX7827,WX8762);
  not NOT_2586(WX7831,WX8762);
  not NOT_2587(WX7833,WX7824);
  not NOT_2588(WX7834,WX7833);
  not NOT_2589(WX7837,WX8761);
  not NOT_2590(WX7841,WX8762);
  not NOT_2591(WX7845,WX8762);
  not NOT_2592(WX7847,WX7838);
  not NOT_2593(WX7848,WX7847);
  not NOT_2594(WX7851,WX8761);
  not NOT_2595(WX7855,WX8762);
  not NOT_2596(WX7859,WX8762);
  not NOT_2597(WX7861,WX7852);
  not NOT_2598(WX7862,WX7861);
  not NOT_2599(WX7865,WX8761);
  not NOT_2600(WX7869,WX8762);
  not NOT_2601(WX7873,WX8762);
  not NOT_2602(WX7875,WX7866);
  not NOT_2603(WX7876,WX7875);
  not NOT_2604(WX7879,WX8761);
  not NOT_2605(WX7883,WX8762);
  not NOT_2606(WX7887,WX8762);
  not NOT_2607(WX7889,WX7880);
  not NOT_2608(WX7890,WX7889);
  not NOT_2609(WX7893,WX8761);
  not NOT_2610(WX7897,WX8762);
  not NOT_2611(WX7901,WX8762);
  not NOT_2612(WX7903,WX7894);
  not NOT_2613(WX7904,WX7903);
  not NOT_2614(WX7907,WX8761);
  not NOT_2615(WX7911,WX8762);
  not NOT_2616(WX7915,WX8762);
  not NOT_2617(WX7917,WX7908);
  not NOT_2618(WX7918,WX7917);
  not NOT_2619(WX7921,WX8761);
  not NOT_2620(WX7925,WX8762);
  not NOT_2621(WX7929,WX8762);
  not NOT_2622(WX7931,WX7922);
  not NOT_2623(WX7932,WX7931);
  not NOT_2624(WX7935,WX8761);
  not NOT_2625(WX7939,WX8762);
  not NOT_2626(WX7943,WX8762);
  not NOT_2627(WX7945,WX7936);
  not NOT_2628(WX7946,WX7945);
  not NOT_2629(WX7949,WX8761);
  not NOT_2630(WX7953,WX8762);
  not NOT_2631(WX7957,WX8762);
  not NOT_2632(WX7959,WX7950);
  not NOT_2633(WX7960,WX7959);
  not NOT_2634(WX7963,WX8761);
  not NOT_2635(WX7967,WX8762);
  not NOT_2636(WX7971,WX8762);
  not NOT_2637(WX7973,WX7964);
  not NOT_2638(WX7974,WX7973);
  not NOT_2639(WX7977,WX8761);
  not NOT_2640(WX7981,WX8762);
  not NOT_2641(WX7985,WX8762);
  not NOT_2642(WX7987,WX7978);
  not NOT_2643(WX7988,WX7987);
  not NOT_2644(WX7991,WX8761);
  not NOT_2645(WX7995,WX8762);
  not NOT_2646(WX7999,WX8762);
  not NOT_2647(WX8001,WX7992);
  not NOT_2648(WX8002,WX8001);
  not NOT_2649(WX8005,WX8761);
  not NOT_2650(WX8009,WX8762);
  not NOT_2651(WX8013,WX8762);
  not NOT_2652(WX8015,WX8006);
  not NOT_2653(WX8016,WX8015);
  not NOT_2654(WX8019,WX8761);
  not NOT_2655(WX8023,WX8762);
  not NOT_2656(WX8027,WX8762);
  not NOT_2657(WX8029,WX8020);
  not NOT_2658(WX8030,WX8029);
  not NOT_2659(WX8033,WX8761);
  not NOT_2660(WX8037,WX8762);
  not NOT_2661(WX8041,WX8762);
  not NOT_2662(WX8043,WX8034);
  not NOT_2663(WX8044,WX8043);
  not NOT_2664(WX8047,WX8761);
  not NOT_2665(WX8051,WX8762);
  not NOT_2666(WX8055,WX8762);
  not NOT_2667(WX8057,WX8048);
  not NOT_2668(WX8058,WX8057);
  not NOT_2669(WX8061,WX8761);
  not NOT_2670(WX8065,WX8762);
  not NOT_2671(WX8069,WX8762);
  not NOT_2672(WX8071,WX8062);
  not NOT_2673(WX8072,WX8071);
  not NOT_2674(WX8075,WX8761);
  not NOT_2675(WX8079,WX8762);
  not NOT_2676(WX8083,WX8762);
  not NOT_2677(WX8085,WX8076);
  not NOT_2678(WX8086,WX8085);
  not NOT_2679(WX8089,WX8761);
  not NOT_2680(WX8093,WX8762);
  not NOT_2681(WX8097,WX8762);
  not NOT_2682(WX8099,WX8090);
  not NOT_2683(WX8100,WX8099);
  not NOT_2684(WX8103,WX8761);
  not NOT_2685(WX8107,WX8762);
  not NOT_2686(WX8111,WX8762);
  not NOT_2687(WX8113,WX8104);
  not NOT_2688(WX8114,WX8113);
  not NOT_2689(WX8117,WX8761);
  not NOT_2690(WX8121,WX8762);
  not NOT_2691(WX8125,WX8762);
  not NOT_2692(WX8127,WX8118);
  not NOT_2693(WX8128,WX8127);
  not NOT_2694(WX8131,WX8761);
  not NOT_2695(WX8135,WX8762);
  not NOT_2696(WX8139,WX8762);
  not NOT_2697(WX8141,WX8132);
  not NOT_2698(WX8142,WX8141);
  not NOT_2699(WX8145,WX8761);
  not NOT_2700(WX8149,WX8762);
  not NOT_2701(WX8153,WX8762);
  not NOT_2702(WX8155,WX8146);
  not NOT_2703(WX8156,WX8155);
  not NOT_2704(WX8159,WX8761);
  not NOT_2705(WX8163,WX8762);
  not NOT_2706(WX8167,WX8762);
  not NOT_2707(WX8169,WX8160);
  not NOT_2708(WX8170,WX8169);
  not NOT_2709(WX8173,WX8761);
  not NOT_2710(WX8177,WX8762);
  not NOT_2711(WX8181,WX8762);
  not NOT_2712(WX8183,WX8174);
  not NOT_2713(WX8184,WX8183);
  not NOT_2714(WX8187,WX8761);
  not NOT_2715(WX8191,WX8762);
  not NOT_2716(WX8195,WX8762);
  not NOT_2717(WX8197,WX8188);
  not NOT_2718(WX8198,WX8197);
  not NOT_2719(WX8201,WX8761);
  not NOT_2720(WX8205,WX8762);
  not NOT_2721(WX8209,WX8762);
  not NOT_2722(WX8211,WX8202);
  not NOT_2723(WX8212,WX8211);
  not NOT_2724(WX8215,WX8761);
  not NOT_2725(WX8219,WX8762);
  not NOT_2726(WX8223,WX8762);
  not NOT_2727(WX8225,WX8216);
  not NOT_2728(WX8226,WX8225);
  not NOT_2729(WX8229,WX8761);
  not NOT_2730(WX8233,WX8762);
  not NOT_2731(WX8237,WX8762);
  not NOT_2732(WX8239,WX8230);
  not NOT_2733(WX8240,WX8239);
  not NOT_2734(WX8241,WX8243);
  not NOT_2735(WX8306,WX8723);
  not NOT_2736(WX8307,WX8725);
  not NOT_2737(WX8308,WX8727);
  not NOT_2738(WX8309,WX8729);
  not NOT_2739(WX8310,WX8731);
  not NOT_2740(WX8311,WX8733);
  not NOT_2741(WX8312,WX8735);
  not NOT_2742(WX8313,WX8737);
  not NOT_2743(WX8314,WX8739);
  not NOT_2744(WX8315,WX8741);
  not NOT_2745(WX8316,WX8743);
  not NOT_2746(WX8317,WX8745);
  not NOT_2747(WX8318,WX8747);
  not NOT_2748(WX8319,WX8749);
  not NOT_2749(WX8320,WX8751);
  not NOT_2750(WX8321,WX8753);
  not NOT_2751(WX8322,WX8691);
  not NOT_2752(WX8323,WX8693);
  not NOT_2753(WX8324,WX8695);
  not NOT_2754(WX8325,WX8697);
  not NOT_2755(WX8326,WX8699);
  not NOT_2756(WX8327,WX8701);
  not NOT_2757(WX8328,WX8703);
  not NOT_2758(WX8329,WX8705);
  not NOT_2759(WX8330,WX8707);
  not NOT_2760(WX8331,WX8709);
  not NOT_2761(WX8332,WX8711);
  not NOT_2762(WX8333,WX8713);
  not NOT_2763(WX8334,WX8715);
  not NOT_2764(WX8335,WX8717);
  not NOT_2765(WX8336,WX8719);
  not NOT_2766(WX8337,WX8721);
  not NOT_2767(WX8338,WX8306);
  not NOT_2768(WX8339,WX8307);
  not NOT_2769(WX8340,WX8308);
  not NOT_2770(WX8341,WX8309);
  not NOT_2771(WX8342,WX8310);
  not NOT_2772(WX8343,WX8311);
  not NOT_2773(WX8344,WX8312);
  not NOT_2774(WX8345,WX8313);
  not NOT_2775(WX8346,WX8314);
  not NOT_2776(WX8347,WX8315);
  not NOT_2777(WX8348,WX8316);
  not NOT_2778(WX8349,WX8317);
  not NOT_2779(WX8350,WX8318);
  not NOT_2780(WX8351,WX8319);
  not NOT_2781(WX8352,WX8320);
  not NOT_2782(WX8353,WX8321);
  not NOT_2783(WX8354,WX8322);
  not NOT_2784(WX8355,WX8323);
  not NOT_2785(WX8356,WX8324);
  not NOT_2786(WX8357,WX8325);
  not NOT_2787(WX8358,WX8326);
  not NOT_2788(WX8359,WX8327);
  not NOT_2789(WX8360,WX8328);
  not NOT_2790(WX8361,WX8329);
  not NOT_2791(WX8362,WX8330);
  not NOT_2792(WX8363,WX8331);
  not NOT_2793(WX8364,WX8332);
  not NOT_2794(WX8365,WX8333);
  not NOT_2795(WX8366,WX8334);
  not NOT_2796(WX8367,WX8335);
  not NOT_2797(WX8368,WX8336);
  not NOT_2798(WX8369,WX8337);
  not NOT_2799(WX8370,WX8595);
  not NOT_2800(WX8371,WX8597);
  not NOT_2801(WX8372,WX8599);
  not NOT_2802(WX8373,WX8601);
  not NOT_2803(WX8374,WX8603);
  not NOT_2804(WX8375,WX8605);
  not NOT_2805(WX8376,WX8607);
  not NOT_2806(WX8377,WX8609);
  not NOT_2807(WX8378,WX8611);
  not NOT_2808(WX8379,WX8613);
  not NOT_2809(WX8380,WX8615);
  not NOT_2810(WX8381,WX8617);
  not NOT_2811(WX8382,WX8619);
  not NOT_2812(WX8383,WX8621);
  not NOT_2813(WX8384,WX8623);
  not NOT_2814(WX8385,WX8625);
  not NOT_2815(WX8386,WX8627);
  not NOT_2816(WX8387,WX8629);
  not NOT_2817(WX8388,WX8631);
  not NOT_2818(WX8389,WX8633);
  not NOT_2819(WX8390,WX8635);
  not NOT_2820(WX8391,WX8637);
  not NOT_2821(WX8392,WX8639);
  not NOT_2822(WX8393,WX8641);
  not NOT_2823(WX8394,WX8643);
  not NOT_2824(WX8395,WX8645);
  not NOT_2825(WX8396,WX8647);
  not NOT_2826(WX8397,WX8649);
  not NOT_2827(WX8398,WX8651);
  not NOT_2828(WX8399,WX8653);
  not NOT_2829(WX8400,WX8655);
  not NOT_2830(WX8401,WX8657);
  not NOT_2831(WX8690,WX8674);
  not NOT_2832(WX8691,WX8690);
  not NOT_2833(WX8692,WX8675);
  not NOT_2834(WX8693,WX8692);
  not NOT_2835(WX8694,WX8676);
  not NOT_2836(WX8695,WX8694);
  not NOT_2837(WX8696,WX8677);
  not NOT_2838(WX8697,WX8696);
  not NOT_2839(WX8698,WX8678);
  not NOT_2840(WX8699,WX8698);
  not NOT_2841(WX8700,WX8679);
  not NOT_2842(WX8701,WX8700);
  not NOT_2843(WX8702,WX8680);
  not NOT_2844(WX8703,WX8702);
  not NOT_2845(WX8704,WX8681);
  not NOT_2846(WX8705,WX8704);
  not NOT_2847(WX8706,WX8682);
  not NOT_2848(WX8707,WX8706);
  not NOT_2849(WX8708,WX8683);
  not NOT_2850(WX8709,WX8708);
  not NOT_2851(WX8710,WX8684);
  not NOT_2852(WX8711,WX8710);
  not NOT_2853(WX8712,WX8685);
  not NOT_2854(WX8713,WX8712);
  not NOT_2855(WX8714,WX8686);
  not NOT_2856(WX8715,WX8714);
  not NOT_2857(WX8716,WX8687);
  not NOT_2858(WX8717,WX8716);
  not NOT_2859(WX8718,WX8688);
  not NOT_2860(WX8719,WX8718);
  not NOT_2861(WX8720,WX8689);
  not NOT_2862(WX8721,WX8720);
  not NOT_2863(WX8722,WX8658);
  not NOT_2864(WX8723,WX8722);
  not NOT_2865(WX8724,WX8659);
  not NOT_2866(WX8725,WX8724);
  not NOT_2867(WX8726,WX8660);
  not NOT_2868(WX8727,WX8726);
  not NOT_2869(WX8728,WX8661);
  not NOT_2870(WX8729,WX8728);
  not NOT_2871(WX8730,WX8662);
  not NOT_2872(WX8731,WX8730);
  not NOT_2873(WX8732,WX8663);
  not NOT_2874(WX8733,WX8732);
  not NOT_2875(WX8734,WX8664);
  not NOT_2876(WX8735,WX8734);
  not NOT_2877(WX8736,WX8665);
  not NOT_2878(WX8737,WX8736);
  not NOT_2879(WX8738,WX8666);
  not NOT_2880(WX8739,WX8738);
  not NOT_2881(WX8740,WX8667);
  not NOT_2882(WX8741,WX8740);
  not NOT_2883(WX8742,WX8668);
  not NOT_2884(WX8743,WX8742);
  not NOT_2885(WX8744,WX8669);
  not NOT_2886(WX8745,WX8744);
  not NOT_2887(WX8746,WX8670);
  not NOT_2888(WX8747,WX8746);
  not NOT_2889(WX8748,WX8671);
  not NOT_2890(WX8749,WX8748);
  not NOT_2891(WX8750,WX8672);
  not NOT_2892(WX8751,WX8750);
  not NOT_2893(WX8752,WX8673);
  not NOT_2894(WX8753,WX8752);
  not NOT_2895(WX8754,TM0);
  not NOT_2896(WX8755,TM0);
  not NOT_2897(WX8756,TM0);
  not NOT_2898(WX8757,TM1);
  not NOT_2899(WX8758,TM1);
  not NOT_2900(WX8759,WX8758);
  not NOT_2901(WX8760,WX8756);
  not NOT_2902(WX8761,WX8757);
  not NOT_2903(WX8762,WX8755);
  not NOT_2904(WX8763,WX8754);
  not NOT_2905(WX8767,WX8763);
  not NOT_2906(WX8769,WX8768);
  not NOT_2907(WX8770,WX8769);
  not NOT_2908(WX8774,WX8763);
  not NOT_2909(WX8776,WX8775);
  not NOT_2910(WX8777,WX8776);
  not NOT_2911(WX8781,WX8763);
  not NOT_2912(WX8783,WX8782);
  not NOT_2913(WX8784,WX8783);
  not NOT_2914(WX8788,WX8763);
  not NOT_2915(WX8790,WX8789);
  not NOT_2916(WX8791,WX8790);
  not NOT_2917(WX8795,WX8763);
  not NOT_2918(WX8797,WX8796);
  not NOT_2919(WX8798,WX8797);
  not NOT_2920(WX8802,WX8763);
  not NOT_2921(WX8804,WX8803);
  not NOT_2922(WX8805,WX8804);
  not NOT_2923(WX8809,WX8763);
  not NOT_2924(WX8811,WX8810);
  not NOT_2925(WX8812,WX8811);
  not NOT_2926(WX8816,WX8763);
  not NOT_2927(WX8818,WX8817);
  not NOT_2928(WX8819,WX8818);
  not NOT_2929(WX8823,WX8763);
  not NOT_2930(WX8825,WX8824);
  not NOT_2931(WX8826,WX8825);
  not NOT_2932(WX8830,WX8763);
  not NOT_2933(WX8832,WX8831);
  not NOT_2934(WX8833,WX8832);
  not NOT_2935(WX8837,WX8763);
  not NOT_2936(WX8839,WX8838);
  not NOT_2937(WX8840,WX8839);
  not NOT_2938(WX8844,WX8763);
  not NOT_2939(WX8846,WX8845);
  not NOT_2940(WX8847,WX8846);
  not NOT_2941(WX8851,WX8763);
  not NOT_2942(WX8853,WX8852);
  not NOT_2943(WX8854,WX8853);
  not NOT_2944(WX8858,WX8763);
  not NOT_2945(WX8860,WX8859);
  not NOT_2946(WX8861,WX8860);
  not NOT_2947(WX8865,WX8763);
  not NOT_2948(WX8867,WX8866);
  not NOT_2949(WX8868,WX8867);
  not NOT_2950(WX8872,WX8763);
  not NOT_2951(WX8874,WX8873);
  not NOT_2952(WX8875,WX8874);
  not NOT_2953(WX8879,WX8763);
  not NOT_2954(WX8881,WX8880);
  not NOT_2955(WX8882,WX8881);
  not NOT_2956(WX8886,WX8763);
  not NOT_2957(WX8888,WX8887);
  not NOT_2958(WX8889,WX8888);
  not NOT_2959(WX8893,WX8763);
  not NOT_2960(WX8895,WX8894);
  not NOT_2961(WX8896,WX8895);
  not NOT_2962(WX8900,WX8763);
  not NOT_2963(WX8902,WX8901);
  not NOT_2964(WX8903,WX8902);
  not NOT_2965(WX8907,WX8763);
  not NOT_2966(WX8909,WX8908);
  not NOT_2967(WX8910,WX8909);
  not NOT_2968(WX8914,WX8763);
  not NOT_2969(WX8916,WX8915);
  not NOT_2970(WX8917,WX8916);
  not NOT_2971(WX8921,WX8763);
  not NOT_2972(WX8923,WX8922);
  not NOT_2973(WX8924,WX8923);
  not NOT_2974(WX8928,WX8763);
  not NOT_2975(WX8930,WX8929);
  not NOT_2976(WX8931,WX8930);
  not NOT_2977(WX8935,WX8763);
  not NOT_2978(WX8937,WX8936);
  not NOT_2979(WX8938,WX8937);
  not NOT_2980(WX8942,WX8763);
  not NOT_2981(WX8944,WX8943);
  not NOT_2982(WX8945,WX8944);
  not NOT_2983(WX8949,WX8763);
  not NOT_2984(WX8951,WX8950);
  not NOT_2985(WX8952,WX8951);
  not NOT_2986(WX8956,WX8763);
  not NOT_2987(WX8958,WX8957);
  not NOT_2988(WX8959,WX8958);
  not NOT_2989(WX8963,WX8763);
  not NOT_2990(WX8965,WX8964);
  not NOT_2991(WX8966,WX8965);
  not NOT_2992(WX8970,WX8763);
  not NOT_2993(WX8972,WX8971);
  not NOT_2994(WX8973,WX8972);
  not NOT_2995(WX8977,WX8763);
  not NOT_2996(WX8979,WX8978);
  not NOT_2997(WX8980,WX8979);
  not NOT_2998(WX8984,WX8763);
  not NOT_2999(WX8986,WX8985);
  not NOT_3000(WX8987,WX8986);
  not NOT_3001(WX8988,RESET);
  not NOT_3002(WX9021,WX8988);
  not NOT_3003(WX9088,WX10054);
  not NOT_3004(WX9092,WX10055);
  not NOT_3005(WX9096,WX10055);
  not NOT_3006(WX9098,WX9089);
  not NOT_3007(WX9099,WX9098);
  not NOT_3008(WX9102,WX10054);
  not NOT_3009(WX9106,WX10055);
  not NOT_3010(WX9110,WX10055);
  not NOT_3011(WX9112,WX9103);
  not NOT_3012(WX9113,WX9112);
  not NOT_3013(WX9116,WX10054);
  not NOT_3014(WX9120,WX10055);
  not NOT_3015(WX9124,WX10055);
  not NOT_3016(WX9126,WX9117);
  not NOT_3017(WX9127,WX9126);
  not NOT_3018(WX9130,WX10054);
  not NOT_3019(WX9134,WX10055);
  not NOT_3020(WX9138,WX10055);
  not NOT_3021(WX9140,WX9131);
  not NOT_3022(WX9141,WX9140);
  not NOT_3023(WX9144,WX10054);
  not NOT_3024(WX9148,WX10055);
  not NOT_3025(WX9152,WX10055);
  not NOT_3026(WX9154,WX9145);
  not NOT_3027(WX9155,WX9154);
  not NOT_3028(WX9158,WX10054);
  not NOT_3029(WX9162,WX10055);
  not NOT_3030(WX9166,WX10055);
  not NOT_3031(WX9168,WX9159);
  not NOT_3032(WX9169,WX9168);
  not NOT_3033(WX9172,WX10054);
  not NOT_3034(WX9176,WX10055);
  not NOT_3035(WX9180,WX10055);
  not NOT_3036(WX9182,WX9173);
  not NOT_3037(WX9183,WX9182);
  not NOT_3038(WX9186,WX10054);
  not NOT_3039(WX9190,WX10055);
  not NOT_3040(WX9194,WX10055);
  not NOT_3041(WX9196,WX9187);
  not NOT_3042(WX9197,WX9196);
  not NOT_3043(WX9200,WX10054);
  not NOT_3044(WX9204,WX10055);
  not NOT_3045(WX9208,WX10055);
  not NOT_3046(WX9210,WX9201);
  not NOT_3047(WX9211,WX9210);
  not NOT_3048(WX9214,WX10054);
  not NOT_3049(WX9218,WX10055);
  not NOT_3050(WX9222,WX10055);
  not NOT_3051(WX9224,WX9215);
  not NOT_3052(WX9225,WX9224);
  not NOT_3053(WX9228,WX10054);
  not NOT_3054(WX9232,WX10055);
  not NOT_3055(WX9236,WX10055);
  not NOT_3056(WX9238,WX9229);
  not NOT_3057(WX9239,WX9238);
  not NOT_3058(WX9242,WX10054);
  not NOT_3059(WX9246,WX10055);
  not NOT_3060(WX9250,WX10055);
  not NOT_3061(WX9252,WX9243);
  not NOT_3062(WX9253,WX9252);
  not NOT_3063(WX9256,WX10054);
  not NOT_3064(WX9260,WX10055);
  not NOT_3065(WX9264,WX10055);
  not NOT_3066(WX9266,WX9257);
  not NOT_3067(WX9267,WX9266);
  not NOT_3068(WX9270,WX10054);
  not NOT_3069(WX9274,WX10055);
  not NOT_3070(WX9278,WX10055);
  not NOT_3071(WX9280,WX9271);
  not NOT_3072(WX9281,WX9280);
  not NOT_3073(WX9284,WX10054);
  not NOT_3074(WX9288,WX10055);
  not NOT_3075(WX9292,WX10055);
  not NOT_3076(WX9294,WX9285);
  not NOT_3077(WX9295,WX9294);
  not NOT_3078(WX9298,WX10054);
  not NOT_3079(WX9302,WX10055);
  not NOT_3080(WX9306,WX10055);
  not NOT_3081(WX9308,WX9299);
  not NOT_3082(WX9309,WX9308);
  not NOT_3083(WX9312,WX10054);
  not NOT_3084(WX9316,WX10055);
  not NOT_3085(WX9320,WX10055);
  not NOT_3086(WX9322,WX9313);
  not NOT_3087(WX9323,WX9322);
  not NOT_3088(WX9326,WX10054);
  not NOT_3089(WX9330,WX10055);
  not NOT_3090(WX9334,WX10055);
  not NOT_3091(WX9336,WX9327);
  not NOT_3092(WX9337,WX9336);
  not NOT_3093(WX9340,WX10054);
  not NOT_3094(WX9344,WX10055);
  not NOT_3095(WX9348,WX10055);
  not NOT_3096(WX9350,WX9341);
  not NOT_3097(WX9351,WX9350);
  not NOT_3098(WX9354,WX10054);
  not NOT_3099(WX9358,WX10055);
  not NOT_3100(WX9362,WX10055);
  not NOT_3101(WX9364,WX9355);
  not NOT_3102(WX9365,WX9364);
  not NOT_3103(WX9368,WX10054);
  not NOT_3104(WX9372,WX10055);
  not NOT_3105(WX9376,WX10055);
  not NOT_3106(WX9378,WX9369);
  not NOT_3107(WX9379,WX9378);
  not NOT_3108(WX9382,WX10054);
  not NOT_3109(WX9386,WX10055);
  not NOT_3110(WX9390,WX10055);
  not NOT_3111(WX9392,WX9383);
  not NOT_3112(WX9393,WX9392);
  not NOT_3113(WX9396,WX10054);
  not NOT_3114(WX9400,WX10055);
  not NOT_3115(WX9404,WX10055);
  not NOT_3116(WX9406,WX9397);
  not NOT_3117(WX9407,WX9406);
  not NOT_3118(WX9410,WX10054);
  not NOT_3119(WX9414,WX10055);
  not NOT_3120(WX9418,WX10055);
  not NOT_3121(WX9420,WX9411);
  not NOT_3122(WX9421,WX9420);
  not NOT_3123(WX9424,WX10054);
  not NOT_3124(WX9428,WX10055);
  not NOT_3125(WX9432,WX10055);
  not NOT_3126(WX9434,WX9425);
  not NOT_3127(WX9435,WX9434);
  not NOT_3128(WX9438,WX10054);
  not NOT_3129(WX9442,WX10055);
  not NOT_3130(WX9446,WX10055);
  not NOT_3131(WX9448,WX9439);
  not NOT_3132(WX9449,WX9448);
  not NOT_3133(WX9452,WX10054);
  not NOT_3134(WX9456,WX10055);
  not NOT_3135(WX9460,WX10055);
  not NOT_3136(WX9462,WX9453);
  not NOT_3137(WX9463,WX9462);
  not NOT_3138(WX9466,WX10054);
  not NOT_3139(WX9470,WX10055);
  not NOT_3140(WX9474,WX10055);
  not NOT_3141(WX9476,WX9467);
  not NOT_3142(WX9477,WX9476);
  not NOT_3143(WX9480,WX10054);
  not NOT_3144(WX9484,WX10055);
  not NOT_3145(WX9488,WX10055);
  not NOT_3146(WX9490,WX9481);
  not NOT_3147(WX9491,WX9490);
  not NOT_3148(WX9494,WX10054);
  not NOT_3149(WX9498,WX10055);
  not NOT_3150(WX9502,WX10055);
  not NOT_3151(WX9504,WX9495);
  not NOT_3152(WX9505,WX9504);
  not NOT_3153(WX9508,WX10054);
  not NOT_3154(WX9512,WX10055);
  not NOT_3155(WX9516,WX10055);
  not NOT_3156(WX9518,WX9509);
  not NOT_3157(WX9519,WX9518);
  not NOT_3158(WX9522,WX10054);
  not NOT_3159(WX9526,WX10055);
  not NOT_3160(WX9530,WX10055);
  not NOT_3161(WX9532,WX9523);
  not NOT_3162(WX9533,WX9532);
  not NOT_3163(WX9534,WX9536);
  not NOT_3164(WX9599,WX10016);
  not NOT_3165(WX9600,WX10018);
  not NOT_3166(WX9601,WX10020);
  not NOT_3167(WX9602,WX10022);
  not NOT_3168(WX9603,WX10024);
  not NOT_3169(WX9604,WX10026);
  not NOT_3170(WX9605,WX10028);
  not NOT_3171(WX9606,WX10030);
  not NOT_3172(WX9607,WX10032);
  not NOT_3173(WX9608,WX10034);
  not NOT_3174(WX9609,WX10036);
  not NOT_3175(WX9610,WX10038);
  not NOT_3176(WX9611,WX10040);
  not NOT_3177(WX9612,WX10042);
  not NOT_3178(WX9613,WX10044);
  not NOT_3179(WX9614,WX10046);
  not NOT_3180(WX9615,WX9984);
  not NOT_3181(WX9616,WX9986);
  not NOT_3182(WX9617,WX9988);
  not NOT_3183(WX9618,WX9990);
  not NOT_3184(WX9619,WX9992);
  not NOT_3185(WX9620,WX9994);
  not NOT_3186(WX9621,WX9996);
  not NOT_3187(WX9622,WX9998);
  not NOT_3188(WX9623,WX10000);
  not NOT_3189(WX9624,WX10002);
  not NOT_3190(WX9625,WX10004);
  not NOT_3191(WX9626,WX10006);
  not NOT_3192(WX9627,WX10008);
  not NOT_3193(WX9628,WX10010);
  not NOT_3194(WX9629,WX10012);
  not NOT_3195(WX9630,WX10014);
  not NOT_3196(WX9631,WX9599);
  not NOT_3197(WX9632,WX9600);
  not NOT_3198(WX9633,WX9601);
  not NOT_3199(WX9634,WX9602);
  not NOT_3200(WX9635,WX9603);
  not NOT_3201(WX9636,WX9604);
  not NOT_3202(WX9637,WX9605);
  not NOT_3203(WX9638,WX9606);
  not NOT_3204(WX9639,WX9607);
  not NOT_3205(WX9640,WX9608);
  not NOT_3206(WX9641,WX9609);
  not NOT_3207(WX9642,WX9610);
  not NOT_3208(WX9643,WX9611);
  not NOT_3209(WX9644,WX9612);
  not NOT_3210(WX9645,WX9613);
  not NOT_3211(WX9646,WX9614);
  not NOT_3212(WX9647,WX9615);
  not NOT_3213(WX9648,WX9616);
  not NOT_3214(WX9649,WX9617);
  not NOT_3215(WX9650,WX9618);
  not NOT_3216(WX9651,WX9619);
  not NOT_3217(WX9652,WX9620);
  not NOT_3218(WX9653,WX9621);
  not NOT_3219(WX9654,WX9622);
  not NOT_3220(WX9655,WX9623);
  not NOT_3221(WX9656,WX9624);
  not NOT_3222(WX9657,WX9625);
  not NOT_3223(WX9658,WX9626);
  not NOT_3224(WX9659,WX9627);
  not NOT_3225(WX9660,WX9628);
  not NOT_3226(WX9661,WX9629);
  not NOT_3227(WX9662,WX9630);
  not NOT_3228(WX9663,WX9888);
  not NOT_3229(WX9664,WX9890);
  not NOT_3230(WX9665,WX9892);
  not NOT_3231(WX9666,WX9894);
  not NOT_3232(WX9667,WX9896);
  not NOT_3233(WX9668,WX9898);
  not NOT_3234(WX9669,WX9900);
  not NOT_3235(WX9670,WX9902);
  not NOT_3236(WX9671,WX9904);
  not NOT_3237(WX9672,WX9906);
  not NOT_3238(WX9673,WX9908);
  not NOT_3239(WX9674,WX9910);
  not NOT_3240(WX9675,WX9912);
  not NOT_3241(WX9676,WX9914);
  not NOT_3242(WX9677,WX9916);
  not NOT_3243(WX9678,WX9918);
  not NOT_3244(WX9679,WX9920);
  not NOT_3245(WX9680,WX9922);
  not NOT_3246(WX9681,WX9924);
  not NOT_3247(WX9682,WX9926);
  not NOT_3248(WX9683,WX9928);
  not NOT_3249(WX9684,WX9930);
  not NOT_3250(WX9685,WX9932);
  not NOT_3251(WX9686,WX9934);
  not NOT_3252(WX9687,WX9936);
  not NOT_3253(WX9688,WX9938);
  not NOT_3254(WX9689,WX9940);
  not NOT_3255(WX9690,WX9942);
  not NOT_3256(WX9691,WX9944);
  not NOT_3257(WX9692,WX9946);
  not NOT_3258(WX9693,WX9948);
  not NOT_3259(WX9694,WX9950);
  not NOT_3260(WX9983,WX9967);
  not NOT_3261(WX9984,WX9983);
  not NOT_3262(WX9985,WX9968);
  not NOT_3263(WX9986,WX9985);
  not NOT_3264(WX9987,WX9969);
  not NOT_3265(WX9988,WX9987);
  not NOT_3266(WX9989,WX9970);
  not NOT_3267(WX9990,WX9989);
  not NOT_3268(WX9991,WX9971);
  not NOT_3269(WX9992,WX9991);
  not NOT_3270(WX9993,WX9972);
  not NOT_3271(WX9994,WX9993);
  not NOT_3272(WX9995,WX9973);
  not NOT_3273(WX9996,WX9995);
  not NOT_3274(WX9997,WX9974);
  not NOT_3275(WX9998,WX9997);
  not NOT_3276(WX9999,WX9975);
  not NOT_3277(WX10000,WX9999);
  not NOT_3278(WX10001,WX9976);
  not NOT_3279(WX10002,WX10001);
  not NOT_3280(WX10003,WX9977);
  not NOT_3281(WX10004,WX10003);
  not NOT_3282(WX10005,WX9978);
  not NOT_3283(WX10006,WX10005);
  not NOT_3284(WX10007,WX9979);
  not NOT_3285(WX10008,WX10007);
  not NOT_3286(WX10009,WX9980);
  not NOT_3287(WX10010,WX10009);
  not NOT_3288(WX10011,WX9981);
  not NOT_3289(WX10012,WX10011);
  not NOT_3290(WX10013,WX9982);
  not NOT_3291(WX10014,WX10013);
  not NOT_3292(WX10015,WX9951);
  not NOT_3293(WX10016,WX10015);
  not NOT_3294(WX10017,WX9952);
  not NOT_3295(WX10018,WX10017);
  not NOT_3296(WX10019,WX9953);
  not NOT_3297(WX10020,WX10019);
  not NOT_3298(WX10021,WX9954);
  not NOT_3299(WX10022,WX10021);
  not NOT_3300(WX10023,WX9955);
  not NOT_3301(WX10024,WX10023);
  not NOT_3302(WX10025,WX9956);
  not NOT_3303(WX10026,WX10025);
  not NOT_3304(WX10027,WX9957);
  not NOT_3305(WX10028,WX10027);
  not NOT_3306(WX10029,WX9958);
  not NOT_3307(WX10030,WX10029);
  not NOT_3308(WX10031,WX9959);
  not NOT_3309(WX10032,WX10031);
  not NOT_3310(WX10033,WX9960);
  not NOT_3311(WX10034,WX10033);
  not NOT_3312(WX10035,WX9961);
  not NOT_3313(WX10036,WX10035);
  not NOT_3314(WX10037,WX9962);
  not NOT_3315(WX10038,WX10037);
  not NOT_3316(WX10039,WX9963);
  not NOT_3317(WX10040,WX10039);
  not NOT_3318(WX10041,WX9964);
  not NOT_3319(WX10042,WX10041);
  not NOT_3320(WX10043,WX9965);
  not NOT_3321(WX10044,WX10043);
  not NOT_3322(WX10045,WX9966);
  not NOT_3323(WX10046,WX10045);
  not NOT_3324(WX10047,TM0);
  not NOT_3325(WX10048,TM0);
  not NOT_3326(WX10049,TM0);
  not NOT_3327(WX10050,TM1);
  not NOT_3328(WX10051,TM1);
  not NOT_3329(WX10052,WX10051);
  not NOT_3330(WX10053,WX10049);
  not NOT_3331(WX10054,WX10050);
  not NOT_3332(WX10055,WX10048);
  not NOT_3333(WX10056,WX10047);
  not NOT_3334(WX10060,WX10056);
  not NOT_3335(WX10062,WX10061);
  not NOT_3336(WX10063,WX10062);
  not NOT_3337(WX10067,WX10056);
  not NOT_3338(WX10069,WX10068);
  not NOT_3339(WX10070,WX10069);
  not NOT_3340(WX10074,WX10056);
  not NOT_3341(WX10076,WX10075);
  not NOT_3342(WX10077,WX10076);
  not NOT_3343(WX10081,WX10056);
  not NOT_3344(WX10083,WX10082);
  not NOT_3345(WX10084,WX10083);
  not NOT_3346(WX10088,WX10056);
  not NOT_3347(WX10090,WX10089);
  not NOT_3348(WX10091,WX10090);
  not NOT_3349(WX10095,WX10056);
  not NOT_3350(WX10097,WX10096);
  not NOT_3351(WX10098,WX10097);
  not NOT_3352(WX10102,WX10056);
  not NOT_3353(WX10104,WX10103);
  not NOT_3354(WX10105,WX10104);
  not NOT_3355(WX10109,WX10056);
  not NOT_3356(WX10111,WX10110);
  not NOT_3357(WX10112,WX10111);
  not NOT_3358(WX10116,WX10056);
  not NOT_3359(WX10118,WX10117);
  not NOT_3360(WX10119,WX10118);
  not NOT_3361(WX10123,WX10056);
  not NOT_3362(WX10125,WX10124);
  not NOT_3363(WX10126,WX10125);
  not NOT_3364(WX10130,WX10056);
  not NOT_3365(WX10132,WX10131);
  not NOT_3366(WX10133,WX10132);
  not NOT_3367(WX10137,WX10056);
  not NOT_3368(WX10139,WX10138);
  not NOT_3369(WX10140,WX10139);
  not NOT_3370(WX10144,WX10056);
  not NOT_3371(WX10146,WX10145);
  not NOT_3372(WX10147,WX10146);
  not NOT_3373(WX10151,WX10056);
  not NOT_3374(WX10153,WX10152);
  not NOT_3375(WX10154,WX10153);
  not NOT_3376(WX10158,WX10056);
  not NOT_3377(WX10160,WX10159);
  not NOT_3378(WX10161,WX10160);
  not NOT_3379(WX10165,WX10056);
  not NOT_3380(WX10167,WX10166);
  not NOT_3381(WX10168,WX10167);
  not NOT_3382(WX10172,WX10056);
  not NOT_3383(WX10174,WX10173);
  not NOT_3384(WX10175,WX10174);
  not NOT_3385(WX10179,WX10056);
  not NOT_3386(WX10181,WX10180);
  not NOT_3387(WX10182,WX10181);
  not NOT_3388(WX10186,WX10056);
  not NOT_3389(WX10188,WX10187);
  not NOT_3390(WX10189,WX10188);
  not NOT_3391(WX10193,WX10056);
  not NOT_3392(WX10195,WX10194);
  not NOT_3393(WX10196,WX10195);
  not NOT_3394(WX10200,WX10056);
  not NOT_3395(WX10202,WX10201);
  not NOT_3396(WX10203,WX10202);
  not NOT_3397(WX10207,WX10056);
  not NOT_3398(WX10209,WX10208);
  not NOT_3399(WX10210,WX10209);
  not NOT_3400(WX10214,WX10056);
  not NOT_3401(WX10216,WX10215);
  not NOT_3402(WX10217,WX10216);
  not NOT_3403(WX10221,WX10056);
  not NOT_3404(WX10223,WX10222);
  not NOT_3405(WX10224,WX10223);
  not NOT_3406(WX10228,WX10056);
  not NOT_3407(WX10230,WX10229);
  not NOT_3408(WX10231,WX10230);
  not NOT_3409(WX10235,WX10056);
  not NOT_3410(WX10237,WX10236);
  not NOT_3411(WX10238,WX10237);
  not NOT_3412(WX10242,WX10056);
  not NOT_3413(WX10244,WX10243);
  not NOT_3414(WX10245,WX10244);
  not NOT_3415(WX10249,WX10056);
  not NOT_3416(WX10251,WX10250);
  not NOT_3417(WX10252,WX10251);
  not NOT_3418(WX10256,WX10056);
  not NOT_3419(WX10258,WX10257);
  not NOT_3420(WX10259,WX10258);
  not NOT_3421(WX10263,WX10056);
  not NOT_3422(WX10265,WX10264);
  not NOT_3423(WX10266,WX10265);
  not NOT_3424(WX10270,WX10056);
  not NOT_3425(WX10272,WX10271);
  not NOT_3426(WX10273,WX10272);
  not NOT_3427(WX10277,WX10056);
  not NOT_3428(WX10279,WX10278);
  not NOT_3429(WX10280,WX10279);
  not NOT_3430(WX10281,RESET);
  not NOT_3431(WX10314,WX10281);
  not NOT_3432(WX10381,WX11347);
  not NOT_3433(WX10385,WX11348);
  not NOT_3434(WX10389,WX11348);
  not NOT_3435(WX10391,WX10382);
  not NOT_3436(WX10392,WX10391);
  not NOT_3437(WX10395,WX11347);
  not NOT_3438(WX10399,WX11348);
  not NOT_3439(WX10403,WX11348);
  not NOT_3440(WX10405,WX10396);
  not NOT_3441(WX10406,WX10405);
  not NOT_3442(WX10409,WX11347);
  not NOT_3443(WX10413,WX11348);
  not NOT_3444(WX10417,WX11348);
  not NOT_3445(WX10419,WX10410);
  not NOT_3446(WX10420,WX10419);
  not NOT_3447(WX10423,WX11347);
  not NOT_3448(WX10427,WX11348);
  not NOT_3449(WX10431,WX11348);
  not NOT_3450(WX10433,WX10424);
  not NOT_3451(WX10434,WX10433);
  not NOT_3452(WX10437,WX11347);
  not NOT_3453(WX10441,WX11348);
  not NOT_3454(WX10445,WX11348);
  not NOT_3455(WX10447,WX10438);
  not NOT_3456(WX10448,WX10447);
  not NOT_3457(WX10451,WX11347);
  not NOT_3458(WX10455,WX11348);
  not NOT_3459(WX10459,WX11348);
  not NOT_3460(WX10461,WX10452);
  not NOT_3461(WX10462,WX10461);
  not NOT_3462(WX10465,WX11347);
  not NOT_3463(WX10469,WX11348);
  not NOT_3464(WX10473,WX11348);
  not NOT_3465(WX10475,WX10466);
  not NOT_3466(WX10476,WX10475);
  not NOT_3467(WX10479,WX11347);
  not NOT_3468(WX10483,WX11348);
  not NOT_3469(WX10487,WX11348);
  not NOT_3470(WX10489,WX10480);
  not NOT_3471(WX10490,WX10489);
  not NOT_3472(WX10493,WX11347);
  not NOT_3473(WX10497,WX11348);
  not NOT_3474(WX10501,WX11348);
  not NOT_3475(WX10503,WX10494);
  not NOT_3476(WX10504,WX10503);
  not NOT_3477(WX10507,WX11347);
  not NOT_3478(WX10511,WX11348);
  not NOT_3479(WX10515,WX11348);
  not NOT_3480(WX10517,WX10508);
  not NOT_3481(WX10518,WX10517);
  not NOT_3482(WX10521,WX11347);
  not NOT_3483(WX10525,WX11348);
  not NOT_3484(WX10529,WX11348);
  not NOT_3485(WX10531,WX10522);
  not NOT_3486(WX10532,WX10531);
  not NOT_3487(WX10535,WX11347);
  not NOT_3488(WX10539,WX11348);
  not NOT_3489(WX10543,WX11348);
  not NOT_3490(WX10545,WX10536);
  not NOT_3491(WX10546,WX10545);
  not NOT_3492(WX10549,WX11347);
  not NOT_3493(WX10553,WX11348);
  not NOT_3494(WX10557,WX11348);
  not NOT_3495(WX10559,WX10550);
  not NOT_3496(WX10560,WX10559);
  not NOT_3497(WX10563,WX11347);
  not NOT_3498(WX10567,WX11348);
  not NOT_3499(WX10571,WX11348);
  not NOT_3500(WX10573,WX10564);
  not NOT_3501(WX10574,WX10573);
  not NOT_3502(WX10577,WX11347);
  not NOT_3503(WX10581,WX11348);
  not NOT_3504(WX10585,WX11348);
  not NOT_3505(WX10587,WX10578);
  not NOT_3506(WX10588,WX10587);
  not NOT_3507(WX10591,WX11347);
  not NOT_3508(WX10595,WX11348);
  not NOT_3509(WX10599,WX11348);
  not NOT_3510(WX10601,WX10592);
  not NOT_3511(WX10602,WX10601);
  not NOT_3512(WX10605,WX11347);
  not NOT_3513(WX10609,WX11348);
  not NOT_3514(WX10613,WX11348);
  not NOT_3515(WX10615,WX10606);
  not NOT_3516(WX10616,WX10615);
  not NOT_3517(WX10619,WX11347);
  not NOT_3518(WX10623,WX11348);
  not NOT_3519(WX10627,WX11348);
  not NOT_3520(WX10629,WX10620);
  not NOT_3521(WX10630,WX10629);
  not NOT_3522(WX10633,WX11347);
  not NOT_3523(WX10637,WX11348);
  not NOT_3524(WX10641,WX11348);
  not NOT_3525(WX10643,WX10634);
  not NOT_3526(WX10644,WX10643);
  not NOT_3527(WX10647,WX11347);
  not NOT_3528(WX10651,WX11348);
  not NOT_3529(WX10655,WX11348);
  not NOT_3530(WX10657,WX10648);
  not NOT_3531(WX10658,WX10657);
  not NOT_3532(WX10661,WX11347);
  not NOT_3533(WX10665,WX11348);
  not NOT_3534(WX10669,WX11348);
  not NOT_3535(WX10671,WX10662);
  not NOT_3536(WX10672,WX10671);
  not NOT_3537(WX10675,WX11347);
  not NOT_3538(WX10679,WX11348);
  not NOT_3539(WX10683,WX11348);
  not NOT_3540(WX10685,WX10676);
  not NOT_3541(WX10686,WX10685);
  not NOT_3542(WX10689,WX11347);
  not NOT_3543(WX10693,WX11348);
  not NOT_3544(WX10697,WX11348);
  not NOT_3545(WX10699,WX10690);
  not NOT_3546(WX10700,WX10699);
  not NOT_3547(WX10703,WX11347);
  not NOT_3548(WX10707,WX11348);
  not NOT_3549(WX10711,WX11348);
  not NOT_3550(WX10713,WX10704);
  not NOT_3551(WX10714,WX10713);
  not NOT_3552(WX10717,WX11347);
  not NOT_3553(WX10721,WX11348);
  not NOT_3554(WX10725,WX11348);
  not NOT_3555(WX10727,WX10718);
  not NOT_3556(WX10728,WX10727);
  not NOT_3557(WX10731,WX11347);
  not NOT_3558(WX10735,WX11348);
  not NOT_3559(WX10739,WX11348);
  not NOT_3560(WX10741,WX10732);
  not NOT_3561(WX10742,WX10741);
  not NOT_3562(WX10745,WX11347);
  not NOT_3563(WX10749,WX11348);
  not NOT_3564(WX10753,WX11348);
  not NOT_3565(WX10755,WX10746);
  not NOT_3566(WX10756,WX10755);
  not NOT_3567(WX10759,WX11347);
  not NOT_3568(WX10763,WX11348);
  not NOT_3569(WX10767,WX11348);
  not NOT_3570(WX10769,WX10760);
  not NOT_3571(WX10770,WX10769);
  not NOT_3572(WX10773,WX11347);
  not NOT_3573(WX10777,WX11348);
  not NOT_3574(WX10781,WX11348);
  not NOT_3575(WX10783,WX10774);
  not NOT_3576(WX10784,WX10783);
  not NOT_3577(WX10787,WX11347);
  not NOT_3578(WX10791,WX11348);
  not NOT_3579(WX10795,WX11348);
  not NOT_3580(WX10797,WX10788);
  not NOT_3581(WX10798,WX10797);
  not NOT_3582(WX10801,WX11347);
  not NOT_3583(WX10805,WX11348);
  not NOT_3584(WX10809,WX11348);
  not NOT_3585(WX10811,WX10802);
  not NOT_3586(WX10812,WX10811);
  not NOT_3587(WX10815,WX11347);
  not NOT_3588(WX10819,WX11348);
  not NOT_3589(WX10823,WX11348);
  not NOT_3590(WX10825,WX10816);
  not NOT_3591(WX10826,WX10825);
  not NOT_3592(WX10827,WX10829);
  not NOT_3593(WX10892,WX11309);
  not NOT_3594(WX10893,WX11311);
  not NOT_3595(WX10894,WX11313);
  not NOT_3596(WX10895,WX11315);
  not NOT_3597(WX10896,WX11317);
  not NOT_3598(WX10897,WX11319);
  not NOT_3599(WX10898,WX11321);
  not NOT_3600(WX10899,WX11323);
  not NOT_3601(WX10900,WX11325);
  not NOT_3602(WX10901,WX11327);
  not NOT_3603(WX10902,WX11329);
  not NOT_3604(WX10903,WX11331);
  not NOT_3605(WX10904,WX11333);
  not NOT_3606(WX10905,WX11335);
  not NOT_3607(WX10906,WX11337);
  not NOT_3608(WX10907,WX11339);
  not NOT_3609(WX10908,WX11277);
  not NOT_3610(WX10909,WX11279);
  not NOT_3611(WX10910,WX11281);
  not NOT_3612(WX10911,WX11283);
  not NOT_3613(WX10912,WX11285);
  not NOT_3614(WX10913,WX11287);
  not NOT_3615(WX10914,WX11289);
  not NOT_3616(WX10915,WX11291);
  not NOT_3617(WX10916,WX11293);
  not NOT_3618(WX10917,WX11295);
  not NOT_3619(WX10918,WX11297);
  not NOT_3620(WX10919,WX11299);
  not NOT_3621(WX10920,WX11301);
  not NOT_3622(WX10921,WX11303);
  not NOT_3623(WX10922,WX11305);
  not NOT_3624(WX10923,WX11307);
  not NOT_3625(WX10924,WX10892);
  not NOT_3626(WX10925,WX10893);
  not NOT_3627(WX10926,WX10894);
  not NOT_3628(WX10927,WX10895);
  not NOT_3629(WX10928,WX10896);
  not NOT_3630(WX10929,WX10897);
  not NOT_3631(WX10930,WX10898);
  not NOT_3632(WX10931,WX10899);
  not NOT_3633(WX10932,WX10900);
  not NOT_3634(WX10933,WX10901);
  not NOT_3635(WX10934,WX10902);
  not NOT_3636(WX10935,WX10903);
  not NOT_3637(WX10936,WX10904);
  not NOT_3638(WX10937,WX10905);
  not NOT_3639(WX10938,WX10906);
  not NOT_3640(WX10939,WX10907);
  not NOT_3641(WX10940,WX10908);
  not NOT_3642(WX10941,WX10909);
  not NOT_3643(WX10942,WX10910);
  not NOT_3644(WX10943,WX10911);
  not NOT_3645(WX10944,WX10912);
  not NOT_3646(WX10945,WX10913);
  not NOT_3647(WX10946,WX10914);
  not NOT_3648(WX10947,WX10915);
  not NOT_3649(WX10948,WX10916);
  not NOT_3650(WX10949,WX10917);
  not NOT_3651(WX10950,WX10918);
  not NOT_3652(WX10951,WX10919);
  not NOT_3653(WX10952,WX10920);
  not NOT_3654(WX10953,WX10921);
  not NOT_3655(WX10954,WX10922);
  not NOT_3656(WX10955,WX10923);
  not NOT_3657(WX10956,WX11181);
  not NOT_3658(WX10957,WX11183);
  not NOT_3659(WX10958,WX11185);
  not NOT_3660(WX10959,WX11187);
  not NOT_3661(WX10960,WX11189);
  not NOT_3662(WX10961,WX11191);
  not NOT_3663(WX10962,WX11193);
  not NOT_3664(WX10963,WX11195);
  not NOT_3665(WX10964,WX11197);
  not NOT_3666(WX10965,WX11199);
  not NOT_3667(WX10966,WX11201);
  not NOT_3668(WX10967,WX11203);
  not NOT_3669(WX10968,WX11205);
  not NOT_3670(WX10969,WX11207);
  not NOT_3671(WX10970,WX11209);
  not NOT_3672(WX10971,WX11211);
  not NOT_3673(WX10972,WX11213);
  not NOT_3674(WX10973,WX11215);
  not NOT_3675(WX10974,WX11217);
  not NOT_3676(WX10975,WX11219);
  not NOT_3677(WX10976,WX11221);
  not NOT_3678(WX10977,WX11223);
  not NOT_3679(WX10978,WX11225);
  not NOT_3680(WX10979,WX11227);
  not NOT_3681(WX10980,WX11229);
  not NOT_3682(WX10981,WX11231);
  not NOT_3683(WX10982,WX11233);
  not NOT_3684(WX10983,WX11235);
  not NOT_3685(WX10984,WX11237);
  not NOT_3686(WX10985,WX11239);
  not NOT_3687(WX10986,WX11241);
  not NOT_3688(WX10987,WX11243);
  not NOT_3689(WX11276,WX11260);
  not NOT_3690(WX11277,WX11276);
  not NOT_3691(WX11278,WX11261);
  not NOT_3692(WX11279,WX11278);
  not NOT_3693(WX11280,WX11262);
  not NOT_3694(WX11281,WX11280);
  not NOT_3695(WX11282,WX11263);
  not NOT_3696(WX11283,WX11282);
  not NOT_3697(WX11284,WX11264);
  not NOT_3698(WX11285,WX11284);
  not NOT_3699(WX11286,WX11265);
  not NOT_3700(WX11287,WX11286);
  not NOT_3701(WX11288,WX11266);
  not NOT_3702(WX11289,WX11288);
  not NOT_3703(WX11290,WX11267);
  not NOT_3704(WX11291,WX11290);
  not NOT_3705(WX11292,WX11268);
  not NOT_3706(WX11293,WX11292);
  not NOT_3707(WX11294,WX11269);
  not NOT_3708(WX11295,WX11294);
  not NOT_3709(WX11296,WX11270);
  not NOT_3710(WX11297,WX11296);
  not NOT_3711(WX11298,WX11271);
  not NOT_3712(WX11299,WX11298);
  not NOT_3713(WX11300,WX11272);
  not NOT_3714(WX11301,WX11300);
  not NOT_3715(WX11302,WX11273);
  not NOT_3716(WX11303,WX11302);
  not NOT_3717(WX11304,WX11274);
  not NOT_3718(WX11305,WX11304);
  not NOT_3719(WX11306,WX11275);
  not NOT_3720(WX11307,WX11306);
  not NOT_3721(WX11308,WX11244);
  not NOT_3722(WX11309,WX11308);
  not NOT_3723(WX11310,WX11245);
  not NOT_3724(WX11311,WX11310);
  not NOT_3725(WX11312,WX11246);
  not NOT_3726(WX11313,WX11312);
  not NOT_3727(WX11314,WX11247);
  not NOT_3728(WX11315,WX11314);
  not NOT_3729(WX11316,WX11248);
  not NOT_3730(WX11317,WX11316);
  not NOT_3731(WX11318,WX11249);
  not NOT_3732(WX11319,WX11318);
  not NOT_3733(WX11320,WX11250);
  not NOT_3734(WX11321,WX11320);
  not NOT_3735(WX11322,WX11251);
  not NOT_3736(WX11323,WX11322);
  not NOT_3737(WX11324,WX11252);
  not NOT_3738(WX11325,WX11324);
  not NOT_3739(WX11326,WX11253);
  not NOT_3740(WX11327,WX11326);
  not NOT_3741(WX11328,WX11254);
  not NOT_3742(WX11329,WX11328);
  not NOT_3743(WX11330,WX11255);
  not NOT_3744(WX11331,WX11330);
  not NOT_3745(WX11332,WX11256);
  not NOT_3746(WX11333,WX11332);
  not NOT_3747(WX11334,WX11257);
  not NOT_3748(WX11335,WX11334);
  not NOT_3749(WX11336,WX11258);
  not NOT_3750(WX11337,WX11336);
  not NOT_3751(WX11338,WX11259);
  not NOT_3752(WX11339,WX11338);
  not NOT_3753(WX11340,TM0);
  not NOT_3754(WX11341,TM0);
  not NOT_3755(WX11342,TM0);
  not NOT_3756(WX11343,TM1);
  not NOT_3757(WX11344,TM1);
  not NOT_3758(WX11345,WX11344);
  not NOT_3759(WX11346,WX11342);
  not NOT_3760(WX11347,WX11343);
  not NOT_3761(WX11348,WX11341);
  not NOT_3762(WX11349,WX11340);
  not NOT_3763(WX11353,WX11349);
  not NOT_3764(WX11355,WX11354);
  not NOT_3765(WX11356,WX11355);
  not NOT_3766(WX11360,WX11349);
  not NOT_3767(WX11362,WX11361);
  not NOT_3768(WX11363,WX11362);
  not NOT_3769(WX11367,WX11349);
  not NOT_3770(WX11369,WX11368);
  not NOT_3771(WX11370,WX11369);
  not NOT_3772(WX11374,WX11349);
  not NOT_3773(WX11376,WX11375);
  not NOT_3774(WX11377,WX11376);
  not NOT_3775(WX11381,WX11349);
  not NOT_3776(WX11383,WX11382);
  not NOT_3777(WX11384,WX11383);
  not NOT_3778(WX11388,WX11349);
  not NOT_3779(WX11390,WX11389);
  not NOT_3780(WX11391,WX11390);
  not NOT_3781(WX11395,WX11349);
  not NOT_3782(WX11397,WX11396);
  not NOT_3783(WX11398,WX11397);
  not NOT_3784(WX11402,WX11349);
  not NOT_3785(WX11404,WX11403);
  not NOT_3786(WX11405,WX11404);
  not NOT_3787(WX11409,WX11349);
  not NOT_3788(WX11411,WX11410);
  not NOT_3789(WX11412,WX11411);
  not NOT_3790(WX11416,WX11349);
  not NOT_3791(WX11418,WX11417);
  not NOT_3792(WX11419,WX11418);
  not NOT_3793(WX11423,WX11349);
  not NOT_3794(WX11425,WX11424);
  not NOT_3795(WX11426,WX11425);
  not NOT_3796(WX11430,WX11349);
  not NOT_3797(WX11432,WX11431);
  not NOT_3798(WX11433,WX11432);
  not NOT_3799(WX11437,WX11349);
  not NOT_3800(WX11439,WX11438);
  not NOT_3801(WX11440,WX11439);
  not NOT_3802(WX11444,WX11349);
  not NOT_3803(WX11446,WX11445);
  not NOT_3804(WX11447,WX11446);
  not NOT_3805(WX11451,WX11349);
  not NOT_3806(WX11453,WX11452);
  not NOT_3807(WX11454,WX11453);
  not NOT_3808(WX11458,WX11349);
  not NOT_3809(WX11460,WX11459);
  not NOT_3810(WX11461,WX11460);
  not NOT_3811(WX11465,WX11349);
  not NOT_3812(WX11467,WX11466);
  not NOT_3813(WX11468,WX11467);
  not NOT_3814(WX11472,WX11349);
  not NOT_3815(WX11474,WX11473);
  not NOT_3816(WX11475,WX11474);
  not NOT_3817(WX11479,WX11349);
  not NOT_3818(WX11481,WX11480);
  not NOT_3819(WX11482,WX11481);
  not NOT_3820(WX11486,WX11349);
  not NOT_3821(WX11488,WX11487);
  not NOT_3822(WX11489,WX11488);
  not NOT_3823(WX11493,WX11349);
  not NOT_3824(WX11495,WX11494);
  not NOT_3825(WX11496,WX11495);
  not NOT_3826(WX11500,WX11349);
  not NOT_3827(WX11502,WX11501);
  not NOT_3828(WX11503,WX11502);
  not NOT_3829(WX11507,WX11349);
  not NOT_3830(WX11509,WX11508);
  not NOT_3831(WX11510,WX11509);
  not NOT_3832(WX11514,WX11349);
  not NOT_3833(WX11516,WX11515);
  not NOT_3834(WX11517,WX11516);
  not NOT_3835(WX11521,WX11349);
  not NOT_3836(WX11523,WX11522);
  not NOT_3837(WX11524,WX11523);
  not NOT_3838(WX11528,WX11349);
  not NOT_3839(WX11530,WX11529);
  not NOT_3840(WX11531,WX11530);
  not NOT_3841(WX11535,WX11349);
  not NOT_3842(WX11537,WX11536);
  not NOT_3843(WX11538,WX11537);
  not NOT_3844(WX11542,WX11349);
  not NOT_3845(WX11544,WX11543);
  not NOT_3846(WX11545,WX11544);
  not NOT_3847(WX11549,WX11349);
  not NOT_3848(WX11551,WX11550);
  not NOT_3849(WX11552,WX11551);
  not NOT_3850(WX11556,WX11349);
  not NOT_3851(WX11558,WX11557);
  not NOT_3852(WX11559,WX11558);
  not NOT_3853(WX11563,WX11349);
  not NOT_3854(WX11565,WX11564);
  not NOT_3855(WX11566,WX11565);
  not NOT_3856(WX11570,WX11349);
  not NOT_3857(WX11572,WX11571);
  not NOT_3858(WX11573,WX11572);
  not NOT_3859(WX11574,RESET);
  not NOT_3860(WX11607,WX11574);
  and AND2_0(WX35,WX46,WX1003);
  and AND2_1(WX36,WX42,WX37);
  and AND2_2(WX39,CRC_OUT_9_31,WX1004);
  and AND2_3(WX40,WX2305,WX41);
  and AND2_4(WX43,WX485,WX1004);
  and AND2_5(WX44,DATA_9_31,WX45);
  and AND2_6(WX49,WX60,WX1003);
  and AND2_7(WX50,WX56,WX51);
  and AND2_8(WX53,CRC_OUT_9_30,WX1004);
  and AND2_9(WX54,WX2312,WX55);
  and AND2_10(WX57,WX487,WX1004);
  and AND2_11(WX58,DATA_9_30,WX59);
  and AND2_12(WX63,WX74,WX1003);
  and AND2_13(WX64,WX70,WX65);
  and AND2_14(WX67,CRC_OUT_9_29,WX1004);
  and AND2_15(WX68,WX2319,WX69);
  and AND2_16(WX71,WX489,WX1004);
  and AND2_17(WX72,DATA_9_29,WX73);
  and AND2_18(WX77,WX88,WX1003);
  and AND2_19(WX78,WX84,WX79);
  and AND2_20(WX81,CRC_OUT_9_28,WX1004);
  and AND2_21(WX82,WX2326,WX83);
  and AND2_22(WX85,WX491,WX1004);
  and AND2_23(WX86,DATA_9_28,WX87);
  and AND2_24(WX91,WX102,WX1003);
  and AND2_25(WX92,WX98,WX93);
  and AND2_26(WX95,CRC_OUT_9_27,WX1004);
  and AND2_27(WX96,WX2333,WX97);
  and AND2_28(WX99,WX493,WX1004);
  and AND2_29(WX100,DATA_9_27,WX101);
  and AND2_30(WX105,WX116,WX1003);
  and AND2_31(WX106,WX112,WX107);
  and AND2_32(WX109,CRC_OUT_9_26,WX1004);
  and AND2_33(WX110,WX2340,WX111);
  and AND2_34(WX113,WX495,WX1004);
  and AND2_35(WX114,DATA_9_26,WX115);
  and AND2_36(WX119,WX130,WX1003);
  and AND2_37(WX120,WX126,WX121);
  and AND2_38(WX123,CRC_OUT_9_25,WX1004);
  and AND2_39(WX124,WX2347,WX125);
  and AND2_40(WX127,WX497,WX1004);
  and AND2_41(WX128,DATA_9_25,WX129);
  and AND2_42(WX133,WX144,WX1003);
  and AND2_43(WX134,WX140,WX135);
  and AND2_44(WX137,CRC_OUT_9_24,WX1004);
  and AND2_45(WX138,WX2354,WX139);
  and AND2_46(WX141,WX499,WX1004);
  and AND2_47(WX142,DATA_9_24,WX143);
  and AND2_48(WX147,WX158,WX1003);
  and AND2_49(WX148,WX154,WX149);
  and AND2_50(WX151,CRC_OUT_9_23,WX1004);
  and AND2_51(WX152,WX2361,WX153);
  and AND2_52(WX155,WX501,WX1004);
  and AND2_53(WX156,DATA_9_23,WX157);
  and AND2_54(WX161,WX172,WX1003);
  and AND2_55(WX162,WX168,WX163);
  and AND2_56(WX165,CRC_OUT_9_22,WX1004);
  and AND2_57(WX166,WX2368,WX167);
  and AND2_58(WX169,WX503,WX1004);
  and AND2_59(WX170,DATA_9_22,WX171);
  and AND2_60(WX175,WX186,WX1003);
  and AND2_61(WX176,WX182,WX177);
  and AND2_62(WX179,CRC_OUT_9_21,WX1004);
  and AND2_63(WX180,WX2375,WX181);
  and AND2_64(WX183,WX505,WX1004);
  and AND2_65(WX184,DATA_9_21,WX185);
  and AND2_66(WX189,WX200,WX1003);
  and AND2_67(WX190,WX196,WX191);
  and AND2_68(WX193,CRC_OUT_9_20,WX1004);
  and AND2_69(WX194,WX2382,WX195);
  and AND2_70(WX197,WX507,WX1004);
  and AND2_71(WX198,DATA_9_20,WX199);
  and AND2_72(WX203,WX214,WX1003);
  and AND2_73(WX204,WX210,WX205);
  and AND2_74(WX207,CRC_OUT_9_19,WX1004);
  and AND2_75(WX208,WX2389,WX209);
  and AND2_76(WX211,WX509,WX1004);
  and AND2_77(WX212,DATA_9_19,WX213);
  and AND2_78(WX217,WX228,WX1003);
  and AND2_79(WX218,WX224,WX219);
  and AND2_80(WX221,CRC_OUT_9_18,WX1004);
  and AND2_81(WX222,WX2396,WX223);
  and AND2_82(WX225,WX511,WX1004);
  and AND2_83(WX226,DATA_9_18,WX227);
  and AND2_84(WX231,WX242,WX1003);
  and AND2_85(WX232,WX238,WX233);
  and AND2_86(WX235,CRC_OUT_9_17,WX1004);
  and AND2_87(WX236,WX2403,WX237);
  and AND2_88(WX239,WX513,WX1004);
  and AND2_89(WX240,DATA_9_17,WX241);
  and AND2_90(WX245,WX256,WX1003);
  and AND2_91(WX246,WX252,WX247);
  and AND2_92(WX249,CRC_OUT_9_16,WX1004);
  and AND2_93(WX250,WX2410,WX251);
  and AND2_94(WX253,WX515,WX1004);
  and AND2_95(WX254,DATA_9_16,WX255);
  and AND2_96(WX259,WX270,WX1003);
  and AND2_97(WX260,WX266,WX261);
  and AND2_98(WX263,CRC_OUT_9_15,WX1004);
  and AND2_99(WX264,WX2417,WX265);
  and AND2_100(WX267,WX517,WX1004);
  and AND2_101(WX268,DATA_9_15,WX269);
  and AND2_102(WX273,WX284,WX1003);
  and AND2_103(WX274,WX280,WX275);
  and AND2_104(WX277,CRC_OUT_9_14,WX1004);
  and AND2_105(WX278,WX2424,WX279);
  and AND2_106(WX281,WX519,WX1004);
  and AND2_107(WX282,DATA_9_14,WX283);
  and AND2_108(WX287,WX298,WX1003);
  and AND2_109(WX288,WX294,WX289);
  and AND2_110(WX291,CRC_OUT_9_13,WX1004);
  and AND2_111(WX292,WX2431,WX293);
  and AND2_112(WX295,WX521,WX1004);
  and AND2_113(WX296,DATA_9_13,WX297);
  and AND2_114(WX301,WX312,WX1003);
  and AND2_115(WX302,WX308,WX303);
  and AND2_116(WX305,CRC_OUT_9_12,WX1004);
  and AND2_117(WX306,WX2438,WX307);
  and AND2_118(WX309,WX523,WX1004);
  and AND2_119(WX310,DATA_9_12,WX311);
  and AND2_120(WX315,WX326,WX1003);
  and AND2_121(WX316,WX322,WX317);
  and AND2_122(WX319,CRC_OUT_9_11,WX1004);
  and AND2_123(WX320,WX2445,WX321);
  and AND2_124(WX323,WX525,WX1004);
  and AND2_125(WX324,DATA_9_11,WX325);
  and AND2_126(WX329,WX340,WX1003);
  and AND2_127(WX330,WX336,WX331);
  and AND2_128(WX333,CRC_OUT_9_10,WX1004);
  and AND2_129(WX334,WX2452,WX335);
  and AND2_130(WX337,WX527,WX1004);
  and AND2_131(WX338,DATA_9_10,WX339);
  and AND2_132(WX343,WX354,WX1003);
  and AND2_133(WX344,WX350,WX345);
  and AND2_134(WX347,CRC_OUT_9_9,WX1004);
  and AND2_135(WX348,WX2459,WX349);
  and AND2_136(WX351,WX529,WX1004);
  and AND2_137(WX352,DATA_9_9,WX353);
  and AND2_138(WX357,WX368,WX1003);
  and AND2_139(WX358,WX364,WX359);
  and AND2_140(WX361,CRC_OUT_9_8,WX1004);
  and AND2_141(WX362,WX2466,WX363);
  and AND2_142(WX365,WX531,WX1004);
  and AND2_143(WX366,DATA_9_8,WX367);
  and AND2_144(WX371,WX382,WX1003);
  and AND2_145(WX372,WX378,WX373);
  and AND2_146(WX375,CRC_OUT_9_7,WX1004);
  and AND2_147(WX376,WX2473,WX377);
  and AND2_148(WX379,WX533,WX1004);
  and AND2_149(WX380,DATA_9_7,WX381);
  and AND2_150(WX385,WX396,WX1003);
  and AND2_151(WX386,WX392,WX387);
  and AND2_152(WX389,CRC_OUT_9_6,WX1004);
  and AND2_153(WX390,WX2480,WX391);
  and AND2_154(WX393,WX535,WX1004);
  and AND2_155(WX394,DATA_9_6,WX395);
  and AND2_156(WX399,WX410,WX1003);
  and AND2_157(WX400,WX406,WX401);
  and AND2_158(WX403,CRC_OUT_9_5,WX1004);
  and AND2_159(WX404,WX2487,WX405);
  and AND2_160(WX407,WX537,WX1004);
  and AND2_161(WX408,DATA_9_5,WX409);
  and AND2_162(WX413,WX424,WX1003);
  and AND2_163(WX414,WX420,WX415);
  and AND2_164(WX417,CRC_OUT_9_4,WX1004);
  and AND2_165(WX418,WX2494,WX419);
  and AND2_166(WX421,WX539,WX1004);
  and AND2_167(WX422,DATA_9_4,WX423);
  and AND2_168(WX427,WX438,WX1003);
  and AND2_169(WX428,WX434,WX429);
  and AND2_170(WX431,CRC_OUT_9_3,WX1004);
  and AND2_171(WX432,WX2501,WX433);
  and AND2_172(WX435,WX541,WX1004);
  and AND2_173(WX436,DATA_9_3,WX437);
  and AND2_174(WX441,WX452,WX1003);
  and AND2_175(WX442,WX448,WX443);
  and AND2_176(WX445,CRC_OUT_9_2,WX1004);
  and AND2_177(WX446,WX2508,WX447);
  and AND2_178(WX449,WX543,WX1004);
  and AND2_179(WX450,DATA_9_2,WX451);
  and AND2_180(WX455,WX466,WX1003);
  and AND2_181(WX456,WX462,WX457);
  and AND2_182(WX459,CRC_OUT_9_1,WX1004);
  and AND2_183(WX460,WX2515,WX461);
  and AND2_184(WX463,WX545,WX1004);
  and AND2_185(WX464,DATA_9_1,WX465);
  and AND2_186(WX469,WX480,WX1003);
  and AND2_187(WX470,WX476,WX471);
  and AND2_188(WX473,CRC_OUT_9_0,WX1004);
  and AND2_189(WX474,WX2522,WX475);
  and AND2_190(WX477,WX547,WX1004);
  and AND2_191(WX478,DATA_9_0,WX479);
  and AND2_192(WX484,WX487,RESET);
  and AND2_193(WX486,WX489,RESET);
  and AND2_194(WX488,WX491,RESET);
  and AND2_195(WX490,WX493,RESET);
  and AND2_196(WX492,WX495,RESET);
  and AND2_197(WX494,WX497,RESET);
  and AND2_198(WX496,WX499,RESET);
  and AND2_199(WX498,WX501,RESET);
  and AND2_200(WX500,WX503,RESET);
  and AND2_201(WX502,WX505,RESET);
  and AND2_202(WX504,WX507,RESET);
  and AND2_203(WX506,WX509,RESET);
  and AND2_204(WX508,WX511,RESET);
  and AND2_205(WX510,WX513,RESET);
  and AND2_206(WX512,WX515,RESET);
  and AND2_207(WX514,WX517,RESET);
  and AND2_208(WX516,WX519,RESET);
  and AND2_209(WX518,WX521,RESET);
  and AND2_210(WX520,WX523,RESET);
  and AND2_211(WX522,WX525,RESET);
  and AND2_212(WX524,WX527,RESET);
  and AND2_213(WX526,WX529,RESET);
  and AND2_214(WX528,WX531,RESET);
  and AND2_215(WX530,WX533,RESET);
  and AND2_216(WX532,WX535,RESET);
  and AND2_217(WX534,WX537,RESET);
  and AND2_218(WX536,WX539,RESET);
  and AND2_219(WX538,WX541,RESET);
  and AND2_220(WX540,WX543,RESET);
  and AND2_221(WX542,WX545,RESET);
  and AND2_222(WX544,WX547,RESET);
  and AND2_223(WX546,WX483,RESET);
  and AND2_224(WX644,WX48,RESET);
  and AND2_225(WX646,WX62,RESET);
  and AND2_226(WX648,WX76,RESET);
  and AND2_227(WX650,WX90,RESET);
  and AND2_228(WX652,WX104,RESET);
  and AND2_229(WX654,WX118,RESET);
  and AND2_230(WX656,WX132,RESET);
  and AND2_231(WX658,WX146,RESET);
  and AND2_232(WX660,WX160,RESET);
  and AND2_233(WX662,WX174,RESET);
  and AND2_234(WX664,WX188,RESET);
  and AND2_235(WX666,WX202,RESET);
  and AND2_236(WX668,WX216,RESET);
  and AND2_237(WX670,WX230,RESET);
  and AND2_238(WX672,WX244,RESET);
  and AND2_239(WX674,WX258,RESET);
  and AND2_240(WX676,WX272,RESET);
  and AND2_241(WX678,WX286,RESET);
  and AND2_242(WX680,WX300,RESET);
  and AND2_243(WX682,WX314,RESET);
  and AND2_244(WX684,WX328,RESET);
  and AND2_245(WX686,WX342,RESET);
  and AND2_246(WX688,WX356,RESET);
  and AND2_247(WX690,WX370,RESET);
  and AND2_248(WX692,WX384,RESET);
  and AND2_249(WX694,WX398,RESET);
  and AND2_250(WX696,WX412,RESET);
  and AND2_251(WX698,WX426,RESET);
  and AND2_252(WX700,WX440,RESET);
  and AND2_253(WX702,WX454,RESET);
  and AND2_254(WX704,WX468,RESET);
  and AND2_255(WX706,WX482,RESET);
  and AND2_256(WX708,WX645,RESET);
  and AND2_257(WX710,WX647,RESET);
  and AND2_258(WX712,WX649,RESET);
  and AND2_259(WX714,WX651,RESET);
  and AND2_260(WX716,WX653,RESET);
  and AND2_261(WX718,WX655,RESET);
  and AND2_262(WX720,WX657,RESET);
  and AND2_263(WX722,WX659,RESET);
  and AND2_264(WX724,WX661,RESET);
  and AND2_265(WX726,WX663,RESET);
  and AND2_266(WX728,WX665,RESET);
  and AND2_267(WX730,WX667,RESET);
  and AND2_268(WX732,WX669,RESET);
  and AND2_269(WX734,WX671,RESET);
  and AND2_270(WX736,WX673,RESET);
  and AND2_271(WX738,WX675,RESET);
  and AND2_272(WX740,WX677,RESET);
  and AND2_273(WX742,WX679,RESET);
  and AND2_274(WX744,WX681,RESET);
  and AND2_275(WX746,WX683,RESET);
  and AND2_276(WX748,WX685,RESET);
  and AND2_277(WX750,WX687,RESET);
  and AND2_278(WX752,WX689,RESET);
  and AND2_279(WX754,WX691,RESET);
  and AND2_280(WX756,WX693,RESET);
  and AND2_281(WX758,WX695,RESET);
  and AND2_282(WX760,WX697,RESET);
  and AND2_283(WX762,WX699,RESET);
  and AND2_284(WX764,WX701,RESET);
  and AND2_285(WX766,WX703,RESET);
  and AND2_286(WX768,WX705,RESET);
  and AND2_287(WX770,WX707,RESET);
  and AND2_288(WX772,WX709,RESET);
  and AND2_289(WX774,WX711,RESET);
  and AND2_290(WX776,WX713,RESET);
  and AND2_291(WX778,WX715,RESET);
  and AND2_292(WX780,WX717,RESET);
  and AND2_293(WX782,WX719,RESET);
  and AND2_294(WX784,WX721,RESET);
  and AND2_295(WX786,WX723,RESET);
  and AND2_296(WX788,WX725,RESET);
  and AND2_297(WX790,WX727,RESET);
  and AND2_298(WX792,WX729,RESET);
  and AND2_299(WX794,WX731,RESET);
  and AND2_300(WX796,WX733,RESET);
  and AND2_301(WX798,WX735,RESET);
  and AND2_302(WX800,WX737,RESET);
  and AND2_303(WX802,WX739,RESET);
  and AND2_304(WX804,WX741,RESET);
  and AND2_305(WX806,WX743,RESET);
  and AND2_306(WX808,WX745,RESET);
  and AND2_307(WX810,WX747,RESET);
  and AND2_308(WX812,WX749,RESET);
  and AND2_309(WX814,WX751,RESET);
  and AND2_310(WX816,WX753,RESET);
  and AND2_311(WX818,WX755,RESET);
  and AND2_312(WX820,WX757,RESET);
  and AND2_313(WX822,WX759,RESET);
  and AND2_314(WX824,WX761,RESET);
  and AND2_315(WX826,WX763,RESET);
  and AND2_316(WX828,WX765,RESET);
  and AND2_317(WX830,WX767,RESET);
  and AND2_318(WX832,WX769,RESET);
  and AND2_319(WX834,WX771,RESET);
  and AND2_320(WX836,WX773,RESET);
  and AND2_321(WX838,WX775,RESET);
  and AND2_322(WX840,WX777,RESET);
  and AND2_323(WX842,WX779,RESET);
  and AND2_324(WX844,WX781,RESET);
  and AND2_325(WX846,WX783,RESET);
  and AND2_326(WX848,WX785,RESET);
  and AND2_327(WX850,WX787,RESET);
  and AND2_328(WX852,WX789,RESET);
  and AND2_329(WX854,WX791,RESET);
  and AND2_330(WX856,WX793,RESET);
  and AND2_331(WX858,WX795,RESET);
  and AND2_332(WX860,WX797,RESET);
  and AND2_333(WX862,WX799,RESET);
  and AND2_334(WX864,WX801,RESET);
  and AND2_335(WX866,WX803,RESET);
  and AND2_336(WX868,WX805,RESET);
  and AND2_337(WX870,WX807,RESET);
  and AND2_338(WX872,WX809,RESET);
  and AND2_339(WX874,WX811,RESET);
  and AND2_340(WX876,WX813,RESET);
  and AND2_341(WX878,WX815,RESET);
  and AND2_342(WX880,WX817,RESET);
  and AND2_343(WX882,WX819,RESET);
  and AND2_344(WX884,WX821,RESET);
  and AND2_345(WX886,WX823,RESET);
  and AND2_346(WX888,WX825,RESET);
  and AND2_347(WX890,WX827,RESET);
  and AND2_348(WX892,WX829,RESET);
  and AND2_349(WX894,WX831,RESET);
  and AND2_350(WX896,WX833,RESET);
  and AND2_351(WX898,WX835,RESET);
  and AND2_352(WX1007,WX1006,WX1005);
  and AND2_353(WX1008,WX580,WX1009);
  and AND2_354(WX1014,WX1013,WX1005);
  and AND2_355(WX1015,WX581,WX1016);
  and AND2_356(WX1021,WX1020,WX1005);
  and AND2_357(WX1022,WX582,WX1023);
  and AND2_358(WX1028,WX1027,WX1005);
  and AND2_359(WX1029,WX583,WX1030);
  and AND2_360(WX1035,WX1034,WX1005);
  and AND2_361(WX1036,WX584,WX1037);
  and AND2_362(WX1042,WX1041,WX1005);
  and AND2_363(WX1043,WX585,WX1044);
  and AND2_364(WX1049,WX1048,WX1005);
  and AND2_365(WX1050,WX586,WX1051);
  and AND2_366(WX1056,WX1055,WX1005);
  and AND2_367(WX1057,WX587,WX1058);
  and AND2_368(WX1063,WX1062,WX1005);
  and AND2_369(WX1064,WX588,WX1065);
  and AND2_370(WX1070,WX1069,WX1005);
  and AND2_371(WX1071,WX589,WX1072);
  and AND2_372(WX1077,WX1076,WX1005);
  and AND2_373(WX1078,WX590,WX1079);
  and AND2_374(WX1084,WX1083,WX1005);
  and AND2_375(WX1085,WX591,WX1086);
  and AND2_376(WX1091,WX1090,WX1005);
  and AND2_377(WX1092,WX592,WX1093);
  and AND2_378(WX1098,WX1097,WX1005);
  and AND2_379(WX1099,WX593,WX1100);
  and AND2_380(WX1105,WX1104,WX1005);
  and AND2_381(WX1106,WX594,WX1107);
  and AND2_382(WX1112,WX1111,WX1005);
  and AND2_383(WX1113,WX595,WX1114);
  and AND2_384(WX1119,WX1118,WX1005);
  and AND2_385(WX1120,WX596,WX1121);
  and AND2_386(WX1126,WX1125,WX1005);
  and AND2_387(WX1127,WX597,WX1128);
  and AND2_388(WX1133,WX1132,WX1005);
  and AND2_389(WX1134,WX598,WX1135);
  and AND2_390(WX1140,WX1139,WX1005);
  and AND2_391(WX1141,WX599,WX1142);
  and AND2_392(WX1147,WX1146,WX1005);
  and AND2_393(WX1148,WX600,WX1149);
  and AND2_394(WX1154,WX1153,WX1005);
  and AND2_395(WX1155,WX601,WX1156);
  and AND2_396(WX1161,WX1160,WX1005);
  and AND2_397(WX1162,WX602,WX1163);
  and AND2_398(WX1168,WX1167,WX1005);
  and AND2_399(WX1169,WX603,WX1170);
  and AND2_400(WX1175,WX1174,WX1005);
  and AND2_401(WX1176,WX604,WX1177);
  and AND2_402(WX1182,WX1181,WX1005);
  and AND2_403(WX1183,WX605,WX1184);
  and AND2_404(WX1189,WX1188,WX1005);
  and AND2_405(WX1190,WX606,WX1191);
  and AND2_406(WX1196,WX1195,WX1005);
  and AND2_407(WX1197,WX607,WX1198);
  and AND2_408(WX1203,WX1202,WX1005);
  and AND2_409(WX1204,WX608,WX1205);
  and AND2_410(WX1210,WX1209,WX1005);
  and AND2_411(WX1211,WX609,WX1212);
  and AND2_412(WX1217,WX1216,WX1005);
  and AND2_413(WX1218,WX610,WX1219);
  and AND2_414(WX1224,WX1223,WX1005);
  and AND2_415(WX1225,WX611,WX1226);
  and AND2_416(WX1264,WX1234,WX1263);
  and AND2_417(WX1266,WX1262,WX1263);
  and AND2_418(WX1268,WX1261,WX1263);
  and AND2_419(WX1270,WX1260,WX1263);
  and AND2_420(WX1272,WX1233,WX1263);
  and AND2_421(WX1274,WX1259,WX1263);
  and AND2_422(WX1276,WX1258,WX1263);
  and AND2_423(WX1278,WX1257,WX1263);
  and AND2_424(WX1280,WX1256,WX1263);
  and AND2_425(WX1282,WX1255,WX1263);
  and AND2_426(WX1284,WX1254,WX1263);
  and AND2_427(WX1286,WX1232,WX1263);
  and AND2_428(WX1288,WX1253,WX1263);
  and AND2_429(WX1290,WX1252,WX1263);
  and AND2_430(WX1292,WX1251,WX1263);
  and AND2_431(WX1294,WX1250,WX1263);
  and AND2_432(WX1296,WX1231,WX1263);
  and AND2_433(WX1298,WX1249,WX1263);
  and AND2_434(WX1300,WX1248,WX1263);
  and AND2_435(WX1302,WX1247,WX1263);
  and AND2_436(WX1304,WX1246,WX1263);
  and AND2_437(WX1306,WX1245,WX1263);
  and AND2_438(WX1308,WX1244,WX1263);
  and AND2_439(WX1310,WX1243,WX1263);
  and AND2_440(WX1312,WX1242,WX1263);
  and AND2_441(WX1314,WX1241,WX1263);
  and AND2_442(WX1316,WX1240,WX1263);
  and AND2_443(WX1318,WX1239,WX1263);
  and AND2_444(WX1320,WX1238,WX1263);
  and AND2_445(WX1322,WX1237,WX1263);
  and AND2_446(WX1324,WX1236,WX1263);
  and AND2_447(WX1326,WX1235,WX1263);
  and AND2_448(WX1328,WX1339,WX2296);
  and AND2_449(WX1329,WX1335,WX1330);
  and AND2_450(WX1332,CRC_OUT_8_31,WX2297);
  and AND2_451(WX1333,WX3598,WX1334);
  and AND2_452(WX1336,WX1778,WX2297);
  and AND2_453(WX1337,WX2305,WX1338);
  and AND2_454(WX1342,WX1353,WX2296);
  and AND2_455(WX1343,WX1349,WX1344);
  and AND2_456(WX1346,CRC_OUT_8_30,WX2297);
  and AND2_457(WX1347,WX3605,WX1348);
  and AND2_458(WX1350,WX1780,WX2297);
  and AND2_459(WX1351,WX2312,WX1352);
  and AND2_460(WX1356,WX1367,WX2296);
  and AND2_461(WX1357,WX1363,WX1358);
  and AND2_462(WX1360,CRC_OUT_8_29,WX2297);
  and AND2_463(WX1361,WX3612,WX1362);
  and AND2_464(WX1364,WX1782,WX2297);
  and AND2_465(WX1365,WX2319,WX1366);
  and AND2_466(WX1370,WX1381,WX2296);
  and AND2_467(WX1371,WX1377,WX1372);
  and AND2_468(WX1374,CRC_OUT_8_28,WX2297);
  and AND2_469(WX1375,WX3619,WX1376);
  and AND2_470(WX1378,WX1784,WX2297);
  and AND2_471(WX1379,WX2326,WX1380);
  and AND2_472(WX1384,WX1395,WX2296);
  and AND2_473(WX1385,WX1391,WX1386);
  and AND2_474(WX1388,CRC_OUT_8_27,WX2297);
  and AND2_475(WX1389,WX3626,WX1390);
  and AND2_476(WX1392,WX1786,WX2297);
  and AND2_477(WX1393,WX2333,WX1394);
  and AND2_478(WX1398,WX1409,WX2296);
  and AND2_479(WX1399,WX1405,WX1400);
  and AND2_480(WX1402,CRC_OUT_8_26,WX2297);
  and AND2_481(WX1403,WX3633,WX1404);
  and AND2_482(WX1406,WX1788,WX2297);
  and AND2_483(WX1407,WX2340,WX1408);
  and AND2_484(WX1412,WX1423,WX2296);
  and AND2_485(WX1413,WX1419,WX1414);
  and AND2_486(WX1416,CRC_OUT_8_25,WX2297);
  and AND2_487(WX1417,WX3640,WX1418);
  and AND2_488(WX1420,WX1790,WX2297);
  and AND2_489(WX1421,WX2347,WX1422);
  and AND2_490(WX1426,WX1437,WX2296);
  and AND2_491(WX1427,WX1433,WX1428);
  and AND2_492(WX1430,CRC_OUT_8_24,WX2297);
  and AND2_493(WX1431,WX3647,WX1432);
  and AND2_494(WX1434,WX1792,WX2297);
  and AND2_495(WX1435,WX2354,WX1436);
  and AND2_496(WX1440,WX1451,WX2296);
  and AND2_497(WX1441,WX1447,WX1442);
  and AND2_498(WX1444,CRC_OUT_8_23,WX2297);
  and AND2_499(WX1445,WX3654,WX1446);
  and AND2_500(WX1448,WX1794,WX2297);
  and AND2_501(WX1449,WX2361,WX1450);
  and AND2_502(WX1454,WX1465,WX2296);
  and AND2_503(WX1455,WX1461,WX1456);
  and AND2_504(WX1458,CRC_OUT_8_22,WX2297);
  and AND2_505(WX1459,WX3661,WX1460);
  and AND2_506(WX1462,WX1796,WX2297);
  and AND2_507(WX1463,WX2368,WX1464);
  and AND2_508(WX1468,WX1479,WX2296);
  and AND2_509(WX1469,WX1475,WX1470);
  and AND2_510(WX1472,CRC_OUT_8_21,WX2297);
  and AND2_511(WX1473,WX3668,WX1474);
  and AND2_512(WX1476,WX1798,WX2297);
  and AND2_513(WX1477,WX2375,WX1478);
  and AND2_514(WX1482,WX1493,WX2296);
  and AND2_515(WX1483,WX1489,WX1484);
  and AND2_516(WX1486,CRC_OUT_8_20,WX2297);
  and AND2_517(WX1487,WX3675,WX1488);
  and AND2_518(WX1490,WX1800,WX2297);
  and AND2_519(WX1491,WX2382,WX1492);
  and AND2_520(WX1496,WX1507,WX2296);
  and AND2_521(WX1497,WX1503,WX1498);
  and AND2_522(WX1500,CRC_OUT_8_19,WX2297);
  and AND2_523(WX1501,WX3682,WX1502);
  and AND2_524(WX1504,WX1802,WX2297);
  and AND2_525(WX1505,WX2389,WX1506);
  and AND2_526(WX1510,WX1521,WX2296);
  and AND2_527(WX1511,WX1517,WX1512);
  and AND2_528(WX1514,CRC_OUT_8_18,WX2297);
  and AND2_529(WX1515,WX3689,WX1516);
  and AND2_530(WX1518,WX1804,WX2297);
  and AND2_531(WX1519,WX2396,WX1520);
  and AND2_532(WX1524,WX1535,WX2296);
  and AND2_533(WX1525,WX1531,WX1526);
  and AND2_534(WX1528,CRC_OUT_8_17,WX2297);
  and AND2_535(WX1529,WX3696,WX1530);
  and AND2_536(WX1532,WX1806,WX2297);
  and AND2_537(WX1533,WX2403,WX1534);
  and AND2_538(WX1538,WX1549,WX2296);
  and AND2_539(WX1539,WX1545,WX1540);
  and AND2_540(WX1542,CRC_OUT_8_16,WX2297);
  and AND2_541(WX1543,WX3703,WX1544);
  and AND2_542(WX1546,WX1808,WX2297);
  and AND2_543(WX1547,WX2410,WX1548);
  and AND2_544(WX1552,WX1563,WX2296);
  and AND2_545(WX1553,WX1559,WX1554);
  and AND2_546(WX1556,CRC_OUT_8_15,WX2297);
  and AND2_547(WX1557,WX3710,WX1558);
  and AND2_548(WX1560,WX1810,WX2297);
  and AND2_549(WX1561,WX2417,WX1562);
  and AND2_550(WX1566,WX1577,WX2296);
  and AND2_551(WX1567,WX1573,WX1568);
  and AND2_552(WX1570,CRC_OUT_8_14,WX2297);
  and AND2_553(WX1571,WX3717,WX1572);
  and AND2_554(WX1574,WX1812,WX2297);
  and AND2_555(WX1575,WX2424,WX1576);
  and AND2_556(WX1580,WX1591,WX2296);
  and AND2_557(WX1581,WX1587,WX1582);
  and AND2_558(WX1584,CRC_OUT_8_13,WX2297);
  and AND2_559(WX1585,WX3724,WX1586);
  and AND2_560(WX1588,WX1814,WX2297);
  and AND2_561(WX1589,WX2431,WX1590);
  and AND2_562(WX1594,WX1605,WX2296);
  and AND2_563(WX1595,WX1601,WX1596);
  and AND2_564(WX1598,CRC_OUT_8_12,WX2297);
  and AND2_565(WX1599,WX3731,WX1600);
  and AND2_566(WX1602,WX1816,WX2297);
  and AND2_567(WX1603,WX2438,WX1604);
  and AND2_568(WX1608,WX1619,WX2296);
  and AND2_569(WX1609,WX1615,WX1610);
  and AND2_570(WX1612,CRC_OUT_8_11,WX2297);
  and AND2_571(WX1613,WX3738,WX1614);
  and AND2_572(WX1616,WX1818,WX2297);
  and AND2_573(WX1617,WX2445,WX1618);
  and AND2_574(WX1622,WX1633,WX2296);
  and AND2_575(WX1623,WX1629,WX1624);
  and AND2_576(WX1626,CRC_OUT_8_10,WX2297);
  and AND2_577(WX1627,WX3745,WX1628);
  and AND2_578(WX1630,WX1820,WX2297);
  and AND2_579(WX1631,WX2452,WX1632);
  and AND2_580(WX1636,WX1647,WX2296);
  and AND2_581(WX1637,WX1643,WX1638);
  and AND2_582(WX1640,CRC_OUT_8_9,WX2297);
  and AND2_583(WX1641,WX3752,WX1642);
  and AND2_584(WX1644,WX1822,WX2297);
  and AND2_585(WX1645,WX2459,WX1646);
  and AND2_586(WX1650,WX1661,WX2296);
  and AND2_587(WX1651,WX1657,WX1652);
  and AND2_588(WX1654,CRC_OUT_8_8,WX2297);
  and AND2_589(WX1655,WX3759,WX1656);
  and AND2_590(WX1658,WX1824,WX2297);
  and AND2_591(WX1659,WX2466,WX1660);
  and AND2_592(WX1664,WX1675,WX2296);
  and AND2_593(WX1665,WX1671,WX1666);
  and AND2_594(WX1668,CRC_OUT_8_7,WX2297);
  and AND2_595(WX1669,WX3766,WX1670);
  and AND2_596(WX1672,WX1826,WX2297);
  and AND2_597(WX1673,WX2473,WX1674);
  and AND2_598(WX1678,WX1689,WX2296);
  and AND2_599(WX1679,WX1685,WX1680);
  and AND2_600(WX1682,CRC_OUT_8_6,WX2297);
  and AND2_601(WX1683,WX3773,WX1684);
  and AND2_602(WX1686,WX1828,WX2297);
  and AND2_603(WX1687,WX2480,WX1688);
  and AND2_604(WX1692,WX1703,WX2296);
  and AND2_605(WX1693,WX1699,WX1694);
  and AND2_606(WX1696,CRC_OUT_8_5,WX2297);
  and AND2_607(WX1697,WX3780,WX1698);
  and AND2_608(WX1700,WX1830,WX2297);
  and AND2_609(WX1701,WX2487,WX1702);
  and AND2_610(WX1706,WX1717,WX2296);
  and AND2_611(WX1707,WX1713,WX1708);
  and AND2_612(WX1710,CRC_OUT_8_4,WX2297);
  and AND2_613(WX1711,WX3787,WX1712);
  and AND2_614(WX1714,WX1832,WX2297);
  and AND2_615(WX1715,WX2494,WX1716);
  and AND2_616(WX1720,WX1731,WX2296);
  and AND2_617(WX1721,WX1727,WX1722);
  and AND2_618(WX1724,CRC_OUT_8_3,WX2297);
  and AND2_619(WX1725,WX3794,WX1726);
  and AND2_620(WX1728,WX1834,WX2297);
  and AND2_621(WX1729,WX2501,WX1730);
  and AND2_622(WX1734,WX1745,WX2296);
  and AND2_623(WX1735,WX1741,WX1736);
  and AND2_624(WX1738,CRC_OUT_8_2,WX2297);
  and AND2_625(WX1739,WX3801,WX1740);
  and AND2_626(WX1742,WX1836,WX2297);
  and AND2_627(WX1743,WX2508,WX1744);
  and AND2_628(WX1748,WX1759,WX2296);
  and AND2_629(WX1749,WX1755,WX1750);
  and AND2_630(WX1752,CRC_OUT_8_1,WX2297);
  and AND2_631(WX1753,WX3808,WX1754);
  and AND2_632(WX1756,WX1838,WX2297);
  and AND2_633(WX1757,WX2515,WX1758);
  and AND2_634(WX1762,WX1773,WX2296);
  and AND2_635(WX1763,WX1769,WX1764);
  and AND2_636(WX1766,CRC_OUT_8_0,WX2297);
  and AND2_637(WX1767,WX3815,WX1768);
  and AND2_638(WX1770,WX1840,WX2297);
  and AND2_639(WX1771,WX2522,WX1772);
  and AND2_640(WX1777,WX1780,RESET);
  and AND2_641(WX1779,WX1782,RESET);
  and AND2_642(WX1781,WX1784,RESET);
  and AND2_643(WX1783,WX1786,RESET);
  and AND2_644(WX1785,WX1788,RESET);
  and AND2_645(WX1787,WX1790,RESET);
  and AND2_646(WX1789,WX1792,RESET);
  and AND2_647(WX1791,WX1794,RESET);
  and AND2_648(WX1793,WX1796,RESET);
  and AND2_649(WX1795,WX1798,RESET);
  and AND2_650(WX1797,WX1800,RESET);
  and AND2_651(WX1799,WX1802,RESET);
  and AND2_652(WX1801,WX1804,RESET);
  and AND2_653(WX1803,WX1806,RESET);
  and AND2_654(WX1805,WX1808,RESET);
  and AND2_655(WX1807,WX1810,RESET);
  and AND2_656(WX1809,WX1812,RESET);
  and AND2_657(WX1811,WX1814,RESET);
  and AND2_658(WX1813,WX1816,RESET);
  and AND2_659(WX1815,WX1818,RESET);
  and AND2_660(WX1817,WX1820,RESET);
  and AND2_661(WX1819,WX1822,RESET);
  and AND2_662(WX1821,WX1824,RESET);
  and AND2_663(WX1823,WX1826,RESET);
  and AND2_664(WX1825,WX1828,RESET);
  and AND2_665(WX1827,WX1830,RESET);
  and AND2_666(WX1829,WX1832,RESET);
  and AND2_667(WX1831,WX1834,RESET);
  and AND2_668(WX1833,WX1836,RESET);
  and AND2_669(WX1835,WX1838,RESET);
  and AND2_670(WX1837,WX1840,RESET);
  and AND2_671(WX1839,WX1776,RESET);
  and AND2_672(WX1937,WX1341,RESET);
  and AND2_673(WX1939,WX1355,RESET);
  and AND2_674(WX1941,WX1369,RESET);
  and AND2_675(WX1943,WX1383,RESET);
  and AND2_676(WX1945,WX1397,RESET);
  and AND2_677(WX1947,WX1411,RESET);
  and AND2_678(WX1949,WX1425,RESET);
  and AND2_679(WX1951,WX1439,RESET);
  and AND2_680(WX1953,WX1453,RESET);
  and AND2_681(WX1955,WX1467,RESET);
  and AND2_682(WX1957,WX1481,RESET);
  and AND2_683(WX1959,WX1495,RESET);
  and AND2_684(WX1961,WX1509,RESET);
  and AND2_685(WX1963,WX1523,RESET);
  and AND2_686(WX1965,WX1537,RESET);
  and AND2_687(WX1967,WX1551,RESET);
  and AND2_688(WX1969,WX1565,RESET);
  and AND2_689(WX1971,WX1579,RESET);
  and AND2_690(WX1973,WX1593,RESET);
  and AND2_691(WX1975,WX1607,RESET);
  and AND2_692(WX1977,WX1621,RESET);
  and AND2_693(WX1979,WX1635,RESET);
  and AND2_694(WX1981,WX1649,RESET);
  and AND2_695(WX1983,WX1663,RESET);
  and AND2_696(WX1985,WX1677,RESET);
  and AND2_697(WX1987,WX1691,RESET);
  and AND2_698(WX1989,WX1705,RESET);
  and AND2_699(WX1991,WX1719,RESET);
  and AND2_700(WX1993,WX1733,RESET);
  and AND2_701(WX1995,WX1747,RESET);
  and AND2_702(WX1997,WX1761,RESET);
  and AND2_703(WX1999,WX1775,RESET);
  and AND2_704(WX2001,WX1938,RESET);
  and AND2_705(WX2003,WX1940,RESET);
  and AND2_706(WX2005,WX1942,RESET);
  and AND2_707(WX2007,WX1944,RESET);
  and AND2_708(WX2009,WX1946,RESET);
  and AND2_709(WX2011,WX1948,RESET);
  and AND2_710(WX2013,WX1950,RESET);
  and AND2_711(WX2015,WX1952,RESET);
  and AND2_712(WX2017,WX1954,RESET);
  and AND2_713(WX2019,WX1956,RESET);
  and AND2_714(WX2021,WX1958,RESET);
  and AND2_715(WX2023,WX1960,RESET);
  and AND2_716(WX2025,WX1962,RESET);
  and AND2_717(WX2027,WX1964,RESET);
  and AND2_718(WX2029,WX1966,RESET);
  and AND2_719(WX2031,WX1968,RESET);
  and AND2_720(WX2033,WX1970,RESET);
  and AND2_721(WX2035,WX1972,RESET);
  and AND2_722(WX2037,WX1974,RESET);
  and AND2_723(WX2039,WX1976,RESET);
  and AND2_724(WX2041,WX1978,RESET);
  and AND2_725(WX2043,WX1980,RESET);
  and AND2_726(WX2045,WX1982,RESET);
  and AND2_727(WX2047,WX1984,RESET);
  and AND2_728(WX2049,WX1986,RESET);
  and AND2_729(WX2051,WX1988,RESET);
  and AND2_730(WX2053,WX1990,RESET);
  and AND2_731(WX2055,WX1992,RESET);
  and AND2_732(WX2057,WX1994,RESET);
  and AND2_733(WX2059,WX1996,RESET);
  and AND2_734(WX2061,WX1998,RESET);
  and AND2_735(WX2063,WX2000,RESET);
  and AND2_736(WX2065,WX2002,RESET);
  and AND2_737(WX2067,WX2004,RESET);
  and AND2_738(WX2069,WX2006,RESET);
  and AND2_739(WX2071,WX2008,RESET);
  and AND2_740(WX2073,WX2010,RESET);
  and AND2_741(WX2075,WX2012,RESET);
  and AND2_742(WX2077,WX2014,RESET);
  and AND2_743(WX2079,WX2016,RESET);
  and AND2_744(WX2081,WX2018,RESET);
  and AND2_745(WX2083,WX2020,RESET);
  and AND2_746(WX2085,WX2022,RESET);
  and AND2_747(WX2087,WX2024,RESET);
  and AND2_748(WX2089,WX2026,RESET);
  and AND2_749(WX2091,WX2028,RESET);
  and AND2_750(WX2093,WX2030,RESET);
  and AND2_751(WX2095,WX2032,RESET);
  and AND2_752(WX2097,WX2034,RESET);
  and AND2_753(WX2099,WX2036,RESET);
  and AND2_754(WX2101,WX2038,RESET);
  and AND2_755(WX2103,WX2040,RESET);
  and AND2_756(WX2105,WX2042,RESET);
  and AND2_757(WX2107,WX2044,RESET);
  and AND2_758(WX2109,WX2046,RESET);
  and AND2_759(WX2111,WX2048,RESET);
  and AND2_760(WX2113,WX2050,RESET);
  and AND2_761(WX2115,WX2052,RESET);
  and AND2_762(WX2117,WX2054,RESET);
  and AND2_763(WX2119,WX2056,RESET);
  and AND2_764(WX2121,WX2058,RESET);
  and AND2_765(WX2123,WX2060,RESET);
  and AND2_766(WX2125,WX2062,RESET);
  and AND2_767(WX2127,WX2064,RESET);
  and AND2_768(WX2129,WX2066,RESET);
  and AND2_769(WX2131,WX2068,RESET);
  and AND2_770(WX2133,WX2070,RESET);
  and AND2_771(WX2135,WX2072,RESET);
  and AND2_772(WX2137,WX2074,RESET);
  and AND2_773(WX2139,WX2076,RESET);
  and AND2_774(WX2141,WX2078,RESET);
  and AND2_775(WX2143,WX2080,RESET);
  and AND2_776(WX2145,WX2082,RESET);
  and AND2_777(WX2147,WX2084,RESET);
  and AND2_778(WX2149,WX2086,RESET);
  and AND2_779(WX2151,WX2088,RESET);
  and AND2_780(WX2153,WX2090,RESET);
  and AND2_781(WX2155,WX2092,RESET);
  and AND2_782(WX2157,WX2094,RESET);
  and AND2_783(WX2159,WX2096,RESET);
  and AND2_784(WX2161,WX2098,RESET);
  and AND2_785(WX2163,WX2100,RESET);
  and AND2_786(WX2165,WX2102,RESET);
  and AND2_787(WX2167,WX2104,RESET);
  and AND2_788(WX2169,WX2106,RESET);
  and AND2_789(WX2171,WX2108,RESET);
  and AND2_790(WX2173,WX2110,RESET);
  and AND2_791(WX2175,WX2112,RESET);
  and AND2_792(WX2177,WX2114,RESET);
  and AND2_793(WX2179,WX2116,RESET);
  and AND2_794(WX2181,WX2118,RESET);
  and AND2_795(WX2183,WX2120,RESET);
  and AND2_796(WX2185,WX2122,RESET);
  and AND2_797(WX2187,WX2124,RESET);
  and AND2_798(WX2189,WX2126,RESET);
  and AND2_799(WX2191,WX2128,RESET);
  and AND2_800(WX2300,WX2299,WX2298);
  and AND2_801(WX2301,WX1873,WX2302);
  and AND2_802(WX2307,WX2306,WX2298);
  and AND2_803(WX2308,WX1874,WX2309);
  and AND2_804(WX2314,WX2313,WX2298);
  and AND2_805(WX2315,WX1875,WX2316);
  and AND2_806(WX2321,WX2320,WX2298);
  and AND2_807(WX2322,WX1876,WX2323);
  and AND2_808(WX2328,WX2327,WX2298);
  and AND2_809(WX2329,WX1877,WX2330);
  and AND2_810(WX2335,WX2334,WX2298);
  and AND2_811(WX2336,WX1878,WX2337);
  and AND2_812(WX2342,WX2341,WX2298);
  and AND2_813(WX2343,WX1879,WX2344);
  and AND2_814(WX2349,WX2348,WX2298);
  and AND2_815(WX2350,WX1880,WX2351);
  and AND2_816(WX2356,WX2355,WX2298);
  and AND2_817(WX2357,WX1881,WX2358);
  and AND2_818(WX2363,WX2362,WX2298);
  and AND2_819(WX2364,WX1882,WX2365);
  and AND2_820(WX2370,WX2369,WX2298);
  and AND2_821(WX2371,WX1883,WX2372);
  and AND2_822(WX2377,WX2376,WX2298);
  and AND2_823(WX2378,WX1884,WX2379);
  and AND2_824(WX2384,WX2383,WX2298);
  and AND2_825(WX2385,WX1885,WX2386);
  and AND2_826(WX2391,WX2390,WX2298);
  and AND2_827(WX2392,WX1886,WX2393);
  and AND2_828(WX2398,WX2397,WX2298);
  and AND2_829(WX2399,WX1887,WX2400);
  and AND2_830(WX2405,WX2404,WX2298);
  and AND2_831(WX2406,WX1888,WX2407);
  and AND2_832(WX2412,WX2411,WX2298);
  and AND2_833(WX2413,WX1889,WX2414);
  and AND2_834(WX2419,WX2418,WX2298);
  and AND2_835(WX2420,WX1890,WX2421);
  and AND2_836(WX2426,WX2425,WX2298);
  and AND2_837(WX2427,WX1891,WX2428);
  and AND2_838(WX2433,WX2432,WX2298);
  and AND2_839(WX2434,WX1892,WX2435);
  and AND2_840(WX2440,WX2439,WX2298);
  and AND2_841(WX2441,WX1893,WX2442);
  and AND2_842(WX2447,WX2446,WX2298);
  and AND2_843(WX2448,WX1894,WX2449);
  and AND2_844(WX2454,WX2453,WX2298);
  and AND2_845(WX2455,WX1895,WX2456);
  and AND2_846(WX2461,WX2460,WX2298);
  and AND2_847(WX2462,WX1896,WX2463);
  and AND2_848(WX2468,WX2467,WX2298);
  and AND2_849(WX2469,WX1897,WX2470);
  and AND2_850(WX2475,WX2474,WX2298);
  and AND2_851(WX2476,WX1898,WX2477);
  and AND2_852(WX2482,WX2481,WX2298);
  and AND2_853(WX2483,WX1899,WX2484);
  and AND2_854(WX2489,WX2488,WX2298);
  and AND2_855(WX2490,WX1900,WX2491);
  and AND2_856(WX2496,WX2495,WX2298);
  and AND2_857(WX2497,WX1901,WX2498);
  and AND2_858(WX2503,WX2502,WX2298);
  and AND2_859(WX2504,WX1902,WX2505);
  and AND2_860(WX2510,WX2509,WX2298);
  and AND2_861(WX2511,WX1903,WX2512);
  and AND2_862(WX2517,WX2516,WX2298);
  and AND2_863(WX2518,WX1904,WX2519);
  and AND2_864(WX2557,WX2527,WX2556);
  and AND2_865(WX2559,WX2555,WX2556);
  and AND2_866(WX2561,WX2554,WX2556);
  and AND2_867(WX2563,WX2553,WX2556);
  and AND2_868(WX2565,WX2526,WX2556);
  and AND2_869(WX2567,WX2552,WX2556);
  and AND2_870(WX2569,WX2551,WX2556);
  and AND2_871(WX2571,WX2550,WX2556);
  and AND2_872(WX2573,WX2549,WX2556);
  and AND2_873(WX2575,WX2548,WX2556);
  and AND2_874(WX2577,WX2547,WX2556);
  and AND2_875(WX2579,WX2525,WX2556);
  and AND2_876(WX2581,WX2546,WX2556);
  and AND2_877(WX2583,WX2545,WX2556);
  and AND2_878(WX2585,WX2544,WX2556);
  and AND2_879(WX2587,WX2543,WX2556);
  and AND2_880(WX2589,WX2524,WX2556);
  and AND2_881(WX2591,WX2542,WX2556);
  and AND2_882(WX2593,WX2541,WX2556);
  and AND2_883(WX2595,WX2540,WX2556);
  and AND2_884(WX2597,WX2539,WX2556);
  and AND2_885(WX2599,WX2538,WX2556);
  and AND2_886(WX2601,WX2537,WX2556);
  and AND2_887(WX2603,WX2536,WX2556);
  and AND2_888(WX2605,WX2535,WX2556);
  and AND2_889(WX2607,WX2534,WX2556);
  and AND2_890(WX2609,WX2533,WX2556);
  and AND2_891(WX2611,WX2532,WX2556);
  and AND2_892(WX2613,WX2531,WX2556);
  and AND2_893(WX2615,WX2530,WX2556);
  and AND2_894(WX2617,WX2529,WX2556);
  and AND2_895(WX2619,WX2528,WX2556);
  and AND2_896(WX2621,WX2632,WX3589);
  and AND2_897(WX2622,WX2628,WX2623);
  and AND2_898(WX2625,CRC_OUT_7_31,WX3590);
  and AND2_899(WX2626,WX4891,WX2627);
  and AND2_900(WX2629,WX3071,WX3590);
  and AND2_901(WX2630,WX3598,WX2631);
  and AND2_902(WX2635,WX2646,WX3589);
  and AND2_903(WX2636,WX2642,WX2637);
  and AND2_904(WX2639,CRC_OUT_7_30,WX3590);
  and AND2_905(WX2640,WX4898,WX2641);
  and AND2_906(WX2643,WX3073,WX3590);
  and AND2_907(WX2644,WX3605,WX2645);
  and AND2_908(WX2649,WX2660,WX3589);
  and AND2_909(WX2650,WX2656,WX2651);
  and AND2_910(WX2653,CRC_OUT_7_29,WX3590);
  and AND2_911(WX2654,WX4905,WX2655);
  and AND2_912(WX2657,WX3075,WX3590);
  and AND2_913(WX2658,WX3612,WX2659);
  and AND2_914(WX2663,WX2674,WX3589);
  and AND2_915(WX2664,WX2670,WX2665);
  and AND2_916(WX2667,CRC_OUT_7_28,WX3590);
  and AND2_917(WX2668,WX4912,WX2669);
  and AND2_918(WX2671,WX3077,WX3590);
  and AND2_919(WX2672,WX3619,WX2673);
  and AND2_920(WX2677,WX2688,WX3589);
  and AND2_921(WX2678,WX2684,WX2679);
  and AND2_922(WX2681,CRC_OUT_7_27,WX3590);
  and AND2_923(WX2682,WX4919,WX2683);
  and AND2_924(WX2685,WX3079,WX3590);
  and AND2_925(WX2686,WX3626,WX2687);
  and AND2_926(WX2691,WX2702,WX3589);
  and AND2_927(WX2692,WX2698,WX2693);
  and AND2_928(WX2695,CRC_OUT_7_26,WX3590);
  and AND2_929(WX2696,WX4926,WX2697);
  and AND2_930(WX2699,WX3081,WX3590);
  and AND2_931(WX2700,WX3633,WX2701);
  and AND2_932(WX2705,WX2716,WX3589);
  and AND2_933(WX2706,WX2712,WX2707);
  and AND2_934(WX2709,CRC_OUT_7_25,WX3590);
  and AND2_935(WX2710,WX4933,WX2711);
  and AND2_936(WX2713,WX3083,WX3590);
  and AND2_937(WX2714,WX3640,WX2715);
  and AND2_938(WX2719,WX2730,WX3589);
  and AND2_939(WX2720,WX2726,WX2721);
  and AND2_940(WX2723,CRC_OUT_7_24,WX3590);
  and AND2_941(WX2724,WX4940,WX2725);
  and AND2_942(WX2727,WX3085,WX3590);
  and AND2_943(WX2728,WX3647,WX2729);
  and AND2_944(WX2733,WX2744,WX3589);
  and AND2_945(WX2734,WX2740,WX2735);
  and AND2_946(WX2737,CRC_OUT_7_23,WX3590);
  and AND2_947(WX2738,WX4947,WX2739);
  and AND2_948(WX2741,WX3087,WX3590);
  and AND2_949(WX2742,WX3654,WX2743);
  and AND2_950(WX2747,WX2758,WX3589);
  and AND2_951(WX2748,WX2754,WX2749);
  and AND2_952(WX2751,CRC_OUT_7_22,WX3590);
  and AND2_953(WX2752,WX4954,WX2753);
  and AND2_954(WX2755,WX3089,WX3590);
  and AND2_955(WX2756,WX3661,WX2757);
  and AND2_956(WX2761,WX2772,WX3589);
  and AND2_957(WX2762,WX2768,WX2763);
  and AND2_958(WX2765,CRC_OUT_7_21,WX3590);
  and AND2_959(WX2766,WX4961,WX2767);
  and AND2_960(WX2769,WX3091,WX3590);
  and AND2_961(WX2770,WX3668,WX2771);
  and AND2_962(WX2775,WX2786,WX3589);
  and AND2_963(WX2776,WX2782,WX2777);
  and AND2_964(WX2779,CRC_OUT_7_20,WX3590);
  and AND2_965(WX2780,WX4968,WX2781);
  and AND2_966(WX2783,WX3093,WX3590);
  and AND2_967(WX2784,WX3675,WX2785);
  and AND2_968(WX2789,WX2800,WX3589);
  and AND2_969(WX2790,WX2796,WX2791);
  and AND2_970(WX2793,CRC_OUT_7_19,WX3590);
  and AND2_971(WX2794,WX4975,WX2795);
  and AND2_972(WX2797,WX3095,WX3590);
  and AND2_973(WX2798,WX3682,WX2799);
  and AND2_974(WX2803,WX2814,WX3589);
  and AND2_975(WX2804,WX2810,WX2805);
  and AND2_976(WX2807,CRC_OUT_7_18,WX3590);
  and AND2_977(WX2808,WX4982,WX2809);
  and AND2_978(WX2811,WX3097,WX3590);
  and AND2_979(WX2812,WX3689,WX2813);
  and AND2_980(WX2817,WX2828,WX3589);
  and AND2_981(WX2818,WX2824,WX2819);
  and AND2_982(WX2821,CRC_OUT_7_17,WX3590);
  and AND2_983(WX2822,WX4989,WX2823);
  and AND2_984(WX2825,WX3099,WX3590);
  and AND2_985(WX2826,WX3696,WX2827);
  and AND2_986(WX2831,WX2842,WX3589);
  and AND2_987(WX2832,WX2838,WX2833);
  and AND2_988(WX2835,CRC_OUT_7_16,WX3590);
  and AND2_989(WX2836,WX4996,WX2837);
  and AND2_990(WX2839,WX3101,WX3590);
  and AND2_991(WX2840,WX3703,WX2841);
  and AND2_992(WX2845,WX2856,WX3589);
  and AND2_993(WX2846,WX2852,WX2847);
  and AND2_994(WX2849,CRC_OUT_7_15,WX3590);
  and AND2_995(WX2850,WX5003,WX2851);
  and AND2_996(WX2853,WX3103,WX3590);
  and AND2_997(WX2854,WX3710,WX2855);
  and AND2_998(WX2859,WX2870,WX3589);
  and AND2_999(WX2860,WX2866,WX2861);
  and AND2_1000(WX2863,CRC_OUT_7_14,WX3590);
  and AND2_1001(WX2864,WX5010,WX2865);
  and AND2_1002(WX2867,WX3105,WX3590);
  and AND2_1003(WX2868,WX3717,WX2869);
  and AND2_1004(WX2873,WX2884,WX3589);
  and AND2_1005(WX2874,WX2880,WX2875);
  and AND2_1006(WX2877,CRC_OUT_7_13,WX3590);
  and AND2_1007(WX2878,WX5017,WX2879);
  and AND2_1008(WX2881,WX3107,WX3590);
  and AND2_1009(WX2882,WX3724,WX2883);
  and AND2_1010(WX2887,WX2898,WX3589);
  and AND2_1011(WX2888,WX2894,WX2889);
  and AND2_1012(WX2891,CRC_OUT_7_12,WX3590);
  and AND2_1013(WX2892,WX5024,WX2893);
  and AND2_1014(WX2895,WX3109,WX3590);
  and AND2_1015(WX2896,WX3731,WX2897);
  and AND2_1016(WX2901,WX2912,WX3589);
  and AND2_1017(WX2902,WX2908,WX2903);
  and AND2_1018(WX2905,CRC_OUT_7_11,WX3590);
  and AND2_1019(WX2906,WX5031,WX2907);
  and AND2_1020(WX2909,WX3111,WX3590);
  and AND2_1021(WX2910,WX3738,WX2911);
  and AND2_1022(WX2915,WX2926,WX3589);
  and AND2_1023(WX2916,WX2922,WX2917);
  and AND2_1024(WX2919,CRC_OUT_7_10,WX3590);
  and AND2_1025(WX2920,WX5038,WX2921);
  and AND2_1026(WX2923,WX3113,WX3590);
  and AND2_1027(WX2924,WX3745,WX2925);
  and AND2_1028(WX2929,WX2940,WX3589);
  and AND2_1029(WX2930,WX2936,WX2931);
  and AND2_1030(WX2933,CRC_OUT_7_9,WX3590);
  and AND2_1031(WX2934,WX5045,WX2935);
  and AND2_1032(WX2937,WX3115,WX3590);
  and AND2_1033(WX2938,WX3752,WX2939);
  and AND2_1034(WX2943,WX2954,WX3589);
  and AND2_1035(WX2944,WX2950,WX2945);
  and AND2_1036(WX2947,CRC_OUT_7_8,WX3590);
  and AND2_1037(WX2948,WX5052,WX2949);
  and AND2_1038(WX2951,WX3117,WX3590);
  and AND2_1039(WX2952,WX3759,WX2953);
  and AND2_1040(WX2957,WX2968,WX3589);
  and AND2_1041(WX2958,WX2964,WX2959);
  and AND2_1042(WX2961,CRC_OUT_7_7,WX3590);
  and AND2_1043(WX2962,WX5059,WX2963);
  and AND2_1044(WX2965,WX3119,WX3590);
  and AND2_1045(WX2966,WX3766,WX2967);
  and AND2_1046(WX2971,WX2982,WX3589);
  and AND2_1047(WX2972,WX2978,WX2973);
  and AND2_1048(WX2975,CRC_OUT_7_6,WX3590);
  and AND2_1049(WX2976,WX5066,WX2977);
  and AND2_1050(WX2979,WX3121,WX3590);
  and AND2_1051(WX2980,WX3773,WX2981);
  and AND2_1052(WX2985,WX2996,WX3589);
  and AND2_1053(WX2986,WX2992,WX2987);
  and AND2_1054(WX2989,CRC_OUT_7_5,WX3590);
  and AND2_1055(WX2990,WX5073,WX2991);
  and AND2_1056(WX2993,WX3123,WX3590);
  and AND2_1057(WX2994,WX3780,WX2995);
  and AND2_1058(WX2999,WX3010,WX3589);
  and AND2_1059(WX3000,WX3006,WX3001);
  and AND2_1060(WX3003,CRC_OUT_7_4,WX3590);
  and AND2_1061(WX3004,WX5080,WX3005);
  and AND2_1062(WX3007,WX3125,WX3590);
  and AND2_1063(WX3008,WX3787,WX3009);
  and AND2_1064(WX3013,WX3024,WX3589);
  and AND2_1065(WX3014,WX3020,WX3015);
  and AND2_1066(WX3017,CRC_OUT_7_3,WX3590);
  and AND2_1067(WX3018,WX5087,WX3019);
  and AND2_1068(WX3021,WX3127,WX3590);
  and AND2_1069(WX3022,WX3794,WX3023);
  and AND2_1070(WX3027,WX3038,WX3589);
  and AND2_1071(WX3028,WX3034,WX3029);
  and AND2_1072(WX3031,CRC_OUT_7_2,WX3590);
  and AND2_1073(WX3032,WX5094,WX3033);
  and AND2_1074(WX3035,WX3129,WX3590);
  and AND2_1075(WX3036,WX3801,WX3037);
  and AND2_1076(WX3041,WX3052,WX3589);
  and AND2_1077(WX3042,WX3048,WX3043);
  and AND2_1078(WX3045,CRC_OUT_7_1,WX3590);
  and AND2_1079(WX3046,WX5101,WX3047);
  and AND2_1080(WX3049,WX3131,WX3590);
  and AND2_1081(WX3050,WX3808,WX3051);
  and AND2_1082(WX3055,WX3066,WX3589);
  and AND2_1083(WX3056,WX3062,WX3057);
  and AND2_1084(WX3059,CRC_OUT_7_0,WX3590);
  and AND2_1085(WX3060,WX5108,WX3061);
  and AND2_1086(WX3063,WX3133,WX3590);
  and AND2_1087(WX3064,WX3815,WX3065);
  and AND2_1088(WX3070,WX3073,RESET);
  and AND2_1089(WX3072,WX3075,RESET);
  and AND2_1090(WX3074,WX3077,RESET);
  and AND2_1091(WX3076,WX3079,RESET);
  and AND2_1092(WX3078,WX3081,RESET);
  and AND2_1093(WX3080,WX3083,RESET);
  and AND2_1094(WX3082,WX3085,RESET);
  and AND2_1095(WX3084,WX3087,RESET);
  and AND2_1096(WX3086,WX3089,RESET);
  and AND2_1097(WX3088,WX3091,RESET);
  and AND2_1098(WX3090,WX3093,RESET);
  and AND2_1099(WX3092,WX3095,RESET);
  and AND2_1100(WX3094,WX3097,RESET);
  and AND2_1101(WX3096,WX3099,RESET);
  and AND2_1102(WX3098,WX3101,RESET);
  and AND2_1103(WX3100,WX3103,RESET);
  and AND2_1104(WX3102,WX3105,RESET);
  and AND2_1105(WX3104,WX3107,RESET);
  and AND2_1106(WX3106,WX3109,RESET);
  and AND2_1107(WX3108,WX3111,RESET);
  and AND2_1108(WX3110,WX3113,RESET);
  and AND2_1109(WX3112,WX3115,RESET);
  and AND2_1110(WX3114,WX3117,RESET);
  and AND2_1111(WX3116,WX3119,RESET);
  and AND2_1112(WX3118,WX3121,RESET);
  and AND2_1113(WX3120,WX3123,RESET);
  and AND2_1114(WX3122,WX3125,RESET);
  and AND2_1115(WX3124,WX3127,RESET);
  and AND2_1116(WX3126,WX3129,RESET);
  and AND2_1117(WX3128,WX3131,RESET);
  and AND2_1118(WX3130,WX3133,RESET);
  and AND2_1119(WX3132,WX3069,RESET);
  and AND2_1120(WX3230,WX2634,RESET);
  and AND2_1121(WX3232,WX2648,RESET);
  and AND2_1122(WX3234,WX2662,RESET);
  and AND2_1123(WX3236,WX2676,RESET);
  and AND2_1124(WX3238,WX2690,RESET);
  and AND2_1125(WX3240,WX2704,RESET);
  and AND2_1126(WX3242,WX2718,RESET);
  and AND2_1127(WX3244,WX2732,RESET);
  and AND2_1128(WX3246,WX2746,RESET);
  and AND2_1129(WX3248,WX2760,RESET);
  and AND2_1130(WX3250,WX2774,RESET);
  and AND2_1131(WX3252,WX2788,RESET);
  and AND2_1132(WX3254,WX2802,RESET);
  and AND2_1133(WX3256,WX2816,RESET);
  and AND2_1134(WX3258,WX2830,RESET);
  and AND2_1135(WX3260,WX2844,RESET);
  and AND2_1136(WX3262,WX2858,RESET);
  and AND2_1137(WX3264,WX2872,RESET);
  and AND2_1138(WX3266,WX2886,RESET);
  and AND2_1139(WX3268,WX2900,RESET);
  and AND2_1140(WX3270,WX2914,RESET);
  and AND2_1141(WX3272,WX2928,RESET);
  and AND2_1142(WX3274,WX2942,RESET);
  and AND2_1143(WX3276,WX2956,RESET);
  and AND2_1144(WX3278,WX2970,RESET);
  and AND2_1145(WX3280,WX2984,RESET);
  and AND2_1146(WX3282,WX2998,RESET);
  and AND2_1147(WX3284,WX3012,RESET);
  and AND2_1148(WX3286,WX3026,RESET);
  and AND2_1149(WX3288,WX3040,RESET);
  and AND2_1150(WX3290,WX3054,RESET);
  and AND2_1151(WX3292,WX3068,RESET);
  and AND2_1152(WX3294,WX3231,RESET);
  and AND2_1153(WX3296,WX3233,RESET);
  and AND2_1154(WX3298,WX3235,RESET);
  and AND2_1155(WX3300,WX3237,RESET);
  and AND2_1156(WX3302,WX3239,RESET);
  and AND2_1157(WX3304,WX3241,RESET);
  and AND2_1158(WX3306,WX3243,RESET);
  and AND2_1159(WX3308,WX3245,RESET);
  and AND2_1160(WX3310,WX3247,RESET);
  and AND2_1161(WX3312,WX3249,RESET);
  and AND2_1162(WX3314,WX3251,RESET);
  and AND2_1163(WX3316,WX3253,RESET);
  and AND2_1164(WX3318,WX3255,RESET);
  and AND2_1165(WX3320,WX3257,RESET);
  and AND2_1166(WX3322,WX3259,RESET);
  and AND2_1167(WX3324,WX3261,RESET);
  and AND2_1168(WX3326,WX3263,RESET);
  and AND2_1169(WX3328,WX3265,RESET);
  and AND2_1170(WX3330,WX3267,RESET);
  and AND2_1171(WX3332,WX3269,RESET);
  and AND2_1172(WX3334,WX3271,RESET);
  and AND2_1173(WX3336,WX3273,RESET);
  and AND2_1174(WX3338,WX3275,RESET);
  and AND2_1175(WX3340,WX3277,RESET);
  and AND2_1176(WX3342,WX3279,RESET);
  and AND2_1177(WX3344,WX3281,RESET);
  and AND2_1178(WX3346,WX3283,RESET);
  and AND2_1179(WX3348,WX3285,RESET);
  and AND2_1180(WX3350,WX3287,RESET);
  and AND2_1181(WX3352,WX3289,RESET);
  and AND2_1182(WX3354,WX3291,RESET);
  and AND2_1183(WX3356,WX3293,RESET);
  and AND2_1184(WX3358,WX3295,RESET);
  and AND2_1185(WX3360,WX3297,RESET);
  and AND2_1186(WX3362,WX3299,RESET);
  and AND2_1187(WX3364,WX3301,RESET);
  and AND2_1188(WX3366,WX3303,RESET);
  and AND2_1189(WX3368,WX3305,RESET);
  and AND2_1190(WX3370,WX3307,RESET);
  and AND2_1191(WX3372,WX3309,RESET);
  and AND2_1192(WX3374,WX3311,RESET);
  and AND2_1193(WX3376,WX3313,RESET);
  and AND2_1194(WX3378,WX3315,RESET);
  and AND2_1195(WX3380,WX3317,RESET);
  and AND2_1196(WX3382,WX3319,RESET);
  and AND2_1197(WX3384,WX3321,RESET);
  and AND2_1198(WX3386,WX3323,RESET);
  and AND2_1199(WX3388,WX3325,RESET);
  and AND2_1200(WX3390,WX3327,RESET);
  and AND2_1201(WX3392,WX3329,RESET);
  and AND2_1202(WX3394,WX3331,RESET);
  and AND2_1203(WX3396,WX3333,RESET);
  and AND2_1204(WX3398,WX3335,RESET);
  and AND2_1205(WX3400,WX3337,RESET);
  and AND2_1206(WX3402,WX3339,RESET);
  and AND2_1207(WX3404,WX3341,RESET);
  and AND2_1208(WX3406,WX3343,RESET);
  and AND2_1209(WX3408,WX3345,RESET);
  and AND2_1210(WX3410,WX3347,RESET);
  and AND2_1211(WX3412,WX3349,RESET);
  and AND2_1212(WX3414,WX3351,RESET);
  and AND2_1213(WX3416,WX3353,RESET);
  and AND2_1214(WX3418,WX3355,RESET);
  and AND2_1215(WX3420,WX3357,RESET);
  and AND2_1216(WX3422,WX3359,RESET);
  and AND2_1217(WX3424,WX3361,RESET);
  and AND2_1218(WX3426,WX3363,RESET);
  and AND2_1219(WX3428,WX3365,RESET);
  and AND2_1220(WX3430,WX3367,RESET);
  and AND2_1221(WX3432,WX3369,RESET);
  and AND2_1222(WX3434,WX3371,RESET);
  and AND2_1223(WX3436,WX3373,RESET);
  and AND2_1224(WX3438,WX3375,RESET);
  and AND2_1225(WX3440,WX3377,RESET);
  and AND2_1226(WX3442,WX3379,RESET);
  and AND2_1227(WX3444,WX3381,RESET);
  and AND2_1228(WX3446,WX3383,RESET);
  and AND2_1229(WX3448,WX3385,RESET);
  and AND2_1230(WX3450,WX3387,RESET);
  and AND2_1231(WX3452,WX3389,RESET);
  and AND2_1232(WX3454,WX3391,RESET);
  and AND2_1233(WX3456,WX3393,RESET);
  and AND2_1234(WX3458,WX3395,RESET);
  and AND2_1235(WX3460,WX3397,RESET);
  and AND2_1236(WX3462,WX3399,RESET);
  and AND2_1237(WX3464,WX3401,RESET);
  and AND2_1238(WX3466,WX3403,RESET);
  and AND2_1239(WX3468,WX3405,RESET);
  and AND2_1240(WX3470,WX3407,RESET);
  and AND2_1241(WX3472,WX3409,RESET);
  and AND2_1242(WX3474,WX3411,RESET);
  and AND2_1243(WX3476,WX3413,RESET);
  and AND2_1244(WX3478,WX3415,RESET);
  and AND2_1245(WX3480,WX3417,RESET);
  and AND2_1246(WX3482,WX3419,RESET);
  and AND2_1247(WX3484,WX3421,RESET);
  and AND2_1248(WX3593,WX3592,WX3591);
  and AND2_1249(WX3594,WX3166,WX3595);
  and AND2_1250(WX3600,WX3599,WX3591);
  and AND2_1251(WX3601,WX3167,WX3602);
  and AND2_1252(WX3607,WX3606,WX3591);
  and AND2_1253(WX3608,WX3168,WX3609);
  and AND2_1254(WX3614,WX3613,WX3591);
  and AND2_1255(WX3615,WX3169,WX3616);
  and AND2_1256(WX3621,WX3620,WX3591);
  and AND2_1257(WX3622,WX3170,WX3623);
  and AND2_1258(WX3628,WX3627,WX3591);
  and AND2_1259(WX3629,WX3171,WX3630);
  and AND2_1260(WX3635,WX3634,WX3591);
  and AND2_1261(WX3636,WX3172,WX3637);
  and AND2_1262(WX3642,WX3641,WX3591);
  and AND2_1263(WX3643,WX3173,WX3644);
  and AND2_1264(WX3649,WX3648,WX3591);
  and AND2_1265(WX3650,WX3174,WX3651);
  and AND2_1266(WX3656,WX3655,WX3591);
  and AND2_1267(WX3657,WX3175,WX3658);
  and AND2_1268(WX3663,WX3662,WX3591);
  and AND2_1269(WX3664,WX3176,WX3665);
  and AND2_1270(WX3670,WX3669,WX3591);
  and AND2_1271(WX3671,WX3177,WX3672);
  and AND2_1272(WX3677,WX3676,WX3591);
  and AND2_1273(WX3678,WX3178,WX3679);
  and AND2_1274(WX3684,WX3683,WX3591);
  and AND2_1275(WX3685,WX3179,WX3686);
  and AND2_1276(WX3691,WX3690,WX3591);
  and AND2_1277(WX3692,WX3180,WX3693);
  and AND2_1278(WX3698,WX3697,WX3591);
  and AND2_1279(WX3699,WX3181,WX3700);
  and AND2_1280(WX3705,WX3704,WX3591);
  and AND2_1281(WX3706,WX3182,WX3707);
  and AND2_1282(WX3712,WX3711,WX3591);
  and AND2_1283(WX3713,WX3183,WX3714);
  and AND2_1284(WX3719,WX3718,WX3591);
  and AND2_1285(WX3720,WX3184,WX3721);
  and AND2_1286(WX3726,WX3725,WX3591);
  and AND2_1287(WX3727,WX3185,WX3728);
  and AND2_1288(WX3733,WX3732,WX3591);
  and AND2_1289(WX3734,WX3186,WX3735);
  and AND2_1290(WX3740,WX3739,WX3591);
  and AND2_1291(WX3741,WX3187,WX3742);
  and AND2_1292(WX3747,WX3746,WX3591);
  and AND2_1293(WX3748,WX3188,WX3749);
  and AND2_1294(WX3754,WX3753,WX3591);
  and AND2_1295(WX3755,WX3189,WX3756);
  and AND2_1296(WX3761,WX3760,WX3591);
  and AND2_1297(WX3762,WX3190,WX3763);
  and AND2_1298(WX3768,WX3767,WX3591);
  and AND2_1299(WX3769,WX3191,WX3770);
  and AND2_1300(WX3775,WX3774,WX3591);
  and AND2_1301(WX3776,WX3192,WX3777);
  and AND2_1302(WX3782,WX3781,WX3591);
  and AND2_1303(WX3783,WX3193,WX3784);
  and AND2_1304(WX3789,WX3788,WX3591);
  and AND2_1305(WX3790,WX3194,WX3791);
  and AND2_1306(WX3796,WX3795,WX3591);
  and AND2_1307(WX3797,WX3195,WX3798);
  and AND2_1308(WX3803,WX3802,WX3591);
  and AND2_1309(WX3804,WX3196,WX3805);
  and AND2_1310(WX3810,WX3809,WX3591);
  and AND2_1311(WX3811,WX3197,WX3812);
  and AND2_1312(WX3850,WX3820,WX3849);
  and AND2_1313(WX3852,WX3848,WX3849);
  and AND2_1314(WX3854,WX3847,WX3849);
  and AND2_1315(WX3856,WX3846,WX3849);
  and AND2_1316(WX3858,WX3819,WX3849);
  and AND2_1317(WX3860,WX3845,WX3849);
  and AND2_1318(WX3862,WX3844,WX3849);
  and AND2_1319(WX3864,WX3843,WX3849);
  and AND2_1320(WX3866,WX3842,WX3849);
  and AND2_1321(WX3868,WX3841,WX3849);
  and AND2_1322(WX3870,WX3840,WX3849);
  and AND2_1323(WX3872,WX3818,WX3849);
  and AND2_1324(WX3874,WX3839,WX3849);
  and AND2_1325(WX3876,WX3838,WX3849);
  and AND2_1326(WX3878,WX3837,WX3849);
  and AND2_1327(WX3880,WX3836,WX3849);
  and AND2_1328(WX3882,WX3817,WX3849);
  and AND2_1329(WX3884,WX3835,WX3849);
  and AND2_1330(WX3886,WX3834,WX3849);
  and AND2_1331(WX3888,WX3833,WX3849);
  and AND2_1332(WX3890,WX3832,WX3849);
  and AND2_1333(WX3892,WX3831,WX3849);
  and AND2_1334(WX3894,WX3830,WX3849);
  and AND2_1335(WX3896,WX3829,WX3849);
  and AND2_1336(WX3898,WX3828,WX3849);
  and AND2_1337(WX3900,WX3827,WX3849);
  and AND2_1338(WX3902,WX3826,WX3849);
  and AND2_1339(WX3904,WX3825,WX3849);
  and AND2_1340(WX3906,WX3824,WX3849);
  and AND2_1341(WX3908,WX3823,WX3849);
  and AND2_1342(WX3910,WX3822,WX3849);
  and AND2_1343(WX3912,WX3821,WX3849);
  and AND2_1344(WX3914,WX3925,WX4882);
  and AND2_1345(WX3915,WX3921,WX3916);
  and AND2_1346(WX3918,CRC_OUT_6_31,WX4883);
  and AND2_1347(WX3919,WX6184,WX3920);
  and AND2_1348(WX3922,WX4364,WX4883);
  and AND2_1349(WX3923,WX4891,WX3924);
  and AND2_1350(WX3928,WX3939,WX4882);
  and AND2_1351(WX3929,WX3935,WX3930);
  and AND2_1352(WX3932,CRC_OUT_6_30,WX4883);
  and AND2_1353(WX3933,WX6191,WX3934);
  and AND2_1354(WX3936,WX4366,WX4883);
  and AND2_1355(WX3937,WX4898,WX3938);
  and AND2_1356(WX3942,WX3953,WX4882);
  and AND2_1357(WX3943,WX3949,WX3944);
  and AND2_1358(WX3946,CRC_OUT_6_29,WX4883);
  and AND2_1359(WX3947,WX6198,WX3948);
  and AND2_1360(WX3950,WX4368,WX4883);
  and AND2_1361(WX3951,WX4905,WX3952);
  and AND2_1362(WX3956,WX3967,WX4882);
  and AND2_1363(WX3957,WX3963,WX3958);
  and AND2_1364(WX3960,CRC_OUT_6_28,WX4883);
  and AND2_1365(WX3961,WX6205,WX3962);
  and AND2_1366(WX3964,WX4370,WX4883);
  and AND2_1367(WX3965,WX4912,WX3966);
  and AND2_1368(WX3970,WX3981,WX4882);
  and AND2_1369(WX3971,WX3977,WX3972);
  and AND2_1370(WX3974,CRC_OUT_6_27,WX4883);
  and AND2_1371(WX3975,WX6212,WX3976);
  and AND2_1372(WX3978,WX4372,WX4883);
  and AND2_1373(WX3979,WX4919,WX3980);
  and AND2_1374(WX3984,WX3995,WX4882);
  and AND2_1375(WX3985,WX3991,WX3986);
  and AND2_1376(WX3988,CRC_OUT_6_26,WX4883);
  and AND2_1377(WX3989,WX6219,WX3990);
  and AND2_1378(WX3992,WX4374,WX4883);
  and AND2_1379(WX3993,WX4926,WX3994);
  and AND2_1380(WX3998,WX4009,WX4882);
  and AND2_1381(WX3999,WX4005,WX4000);
  and AND2_1382(WX4002,CRC_OUT_6_25,WX4883);
  and AND2_1383(WX4003,WX6226,WX4004);
  and AND2_1384(WX4006,WX4376,WX4883);
  and AND2_1385(WX4007,WX4933,WX4008);
  and AND2_1386(WX4012,WX4023,WX4882);
  and AND2_1387(WX4013,WX4019,WX4014);
  and AND2_1388(WX4016,CRC_OUT_6_24,WX4883);
  and AND2_1389(WX4017,WX6233,WX4018);
  and AND2_1390(WX4020,WX4378,WX4883);
  and AND2_1391(WX4021,WX4940,WX4022);
  and AND2_1392(WX4026,WX4037,WX4882);
  and AND2_1393(WX4027,WX4033,WX4028);
  and AND2_1394(WX4030,CRC_OUT_6_23,WX4883);
  and AND2_1395(WX4031,WX6240,WX4032);
  and AND2_1396(WX4034,WX4380,WX4883);
  and AND2_1397(WX4035,WX4947,WX4036);
  and AND2_1398(WX4040,WX4051,WX4882);
  and AND2_1399(WX4041,WX4047,WX4042);
  and AND2_1400(WX4044,CRC_OUT_6_22,WX4883);
  and AND2_1401(WX4045,WX6247,WX4046);
  and AND2_1402(WX4048,WX4382,WX4883);
  and AND2_1403(WX4049,WX4954,WX4050);
  and AND2_1404(WX4054,WX4065,WX4882);
  and AND2_1405(WX4055,WX4061,WX4056);
  and AND2_1406(WX4058,CRC_OUT_6_21,WX4883);
  and AND2_1407(WX4059,WX6254,WX4060);
  and AND2_1408(WX4062,WX4384,WX4883);
  and AND2_1409(WX4063,WX4961,WX4064);
  and AND2_1410(WX4068,WX4079,WX4882);
  and AND2_1411(WX4069,WX4075,WX4070);
  and AND2_1412(WX4072,CRC_OUT_6_20,WX4883);
  and AND2_1413(WX4073,WX6261,WX4074);
  and AND2_1414(WX4076,WX4386,WX4883);
  and AND2_1415(WX4077,WX4968,WX4078);
  and AND2_1416(WX4082,WX4093,WX4882);
  and AND2_1417(WX4083,WX4089,WX4084);
  and AND2_1418(WX4086,CRC_OUT_6_19,WX4883);
  and AND2_1419(WX4087,WX6268,WX4088);
  and AND2_1420(WX4090,WX4388,WX4883);
  and AND2_1421(WX4091,WX4975,WX4092);
  and AND2_1422(WX4096,WX4107,WX4882);
  and AND2_1423(WX4097,WX4103,WX4098);
  and AND2_1424(WX4100,CRC_OUT_6_18,WX4883);
  and AND2_1425(WX4101,WX6275,WX4102);
  and AND2_1426(WX4104,WX4390,WX4883);
  and AND2_1427(WX4105,WX4982,WX4106);
  and AND2_1428(WX4110,WX4121,WX4882);
  and AND2_1429(WX4111,WX4117,WX4112);
  and AND2_1430(WX4114,CRC_OUT_6_17,WX4883);
  and AND2_1431(WX4115,WX6282,WX4116);
  and AND2_1432(WX4118,WX4392,WX4883);
  and AND2_1433(WX4119,WX4989,WX4120);
  and AND2_1434(WX4124,WX4135,WX4882);
  and AND2_1435(WX4125,WX4131,WX4126);
  and AND2_1436(WX4128,CRC_OUT_6_16,WX4883);
  and AND2_1437(WX4129,WX6289,WX4130);
  and AND2_1438(WX4132,WX4394,WX4883);
  and AND2_1439(WX4133,WX4996,WX4134);
  and AND2_1440(WX4138,WX4149,WX4882);
  and AND2_1441(WX4139,WX4145,WX4140);
  and AND2_1442(WX4142,CRC_OUT_6_15,WX4883);
  and AND2_1443(WX4143,WX6296,WX4144);
  and AND2_1444(WX4146,WX4396,WX4883);
  and AND2_1445(WX4147,WX5003,WX4148);
  and AND2_1446(WX4152,WX4163,WX4882);
  and AND2_1447(WX4153,WX4159,WX4154);
  and AND2_1448(WX4156,CRC_OUT_6_14,WX4883);
  and AND2_1449(WX4157,WX6303,WX4158);
  and AND2_1450(WX4160,WX4398,WX4883);
  and AND2_1451(WX4161,WX5010,WX4162);
  and AND2_1452(WX4166,WX4177,WX4882);
  and AND2_1453(WX4167,WX4173,WX4168);
  and AND2_1454(WX4170,CRC_OUT_6_13,WX4883);
  and AND2_1455(WX4171,WX6310,WX4172);
  and AND2_1456(WX4174,WX4400,WX4883);
  and AND2_1457(WX4175,WX5017,WX4176);
  and AND2_1458(WX4180,WX4191,WX4882);
  and AND2_1459(WX4181,WX4187,WX4182);
  and AND2_1460(WX4184,CRC_OUT_6_12,WX4883);
  and AND2_1461(WX4185,WX6317,WX4186);
  and AND2_1462(WX4188,WX4402,WX4883);
  and AND2_1463(WX4189,WX5024,WX4190);
  and AND2_1464(WX4194,WX4205,WX4882);
  and AND2_1465(WX4195,WX4201,WX4196);
  and AND2_1466(WX4198,CRC_OUT_6_11,WX4883);
  and AND2_1467(WX4199,WX6324,WX4200);
  and AND2_1468(WX4202,WX4404,WX4883);
  and AND2_1469(WX4203,WX5031,WX4204);
  and AND2_1470(WX4208,WX4219,WX4882);
  and AND2_1471(WX4209,WX4215,WX4210);
  and AND2_1472(WX4212,CRC_OUT_6_10,WX4883);
  and AND2_1473(WX4213,WX6331,WX4214);
  and AND2_1474(WX4216,WX4406,WX4883);
  and AND2_1475(WX4217,WX5038,WX4218);
  and AND2_1476(WX4222,WX4233,WX4882);
  and AND2_1477(WX4223,WX4229,WX4224);
  and AND2_1478(WX4226,CRC_OUT_6_9,WX4883);
  and AND2_1479(WX4227,WX6338,WX4228);
  and AND2_1480(WX4230,WX4408,WX4883);
  and AND2_1481(WX4231,WX5045,WX4232);
  and AND2_1482(WX4236,WX4247,WX4882);
  and AND2_1483(WX4237,WX4243,WX4238);
  and AND2_1484(WX4240,CRC_OUT_6_8,WX4883);
  and AND2_1485(WX4241,WX6345,WX4242);
  and AND2_1486(WX4244,WX4410,WX4883);
  and AND2_1487(WX4245,WX5052,WX4246);
  and AND2_1488(WX4250,WX4261,WX4882);
  and AND2_1489(WX4251,WX4257,WX4252);
  and AND2_1490(WX4254,CRC_OUT_6_7,WX4883);
  and AND2_1491(WX4255,WX6352,WX4256);
  and AND2_1492(WX4258,WX4412,WX4883);
  and AND2_1493(WX4259,WX5059,WX4260);
  and AND2_1494(WX4264,WX4275,WX4882);
  and AND2_1495(WX4265,WX4271,WX4266);
  and AND2_1496(WX4268,CRC_OUT_6_6,WX4883);
  and AND2_1497(WX4269,WX6359,WX4270);
  and AND2_1498(WX4272,WX4414,WX4883);
  and AND2_1499(WX4273,WX5066,WX4274);
  and AND2_1500(WX4278,WX4289,WX4882);
  and AND2_1501(WX4279,WX4285,WX4280);
  and AND2_1502(WX4282,CRC_OUT_6_5,WX4883);
  and AND2_1503(WX4283,WX6366,WX4284);
  and AND2_1504(WX4286,WX4416,WX4883);
  and AND2_1505(WX4287,WX5073,WX4288);
  and AND2_1506(WX4292,WX4303,WX4882);
  and AND2_1507(WX4293,WX4299,WX4294);
  and AND2_1508(WX4296,CRC_OUT_6_4,WX4883);
  and AND2_1509(WX4297,WX6373,WX4298);
  and AND2_1510(WX4300,WX4418,WX4883);
  and AND2_1511(WX4301,WX5080,WX4302);
  and AND2_1512(WX4306,WX4317,WX4882);
  and AND2_1513(WX4307,WX4313,WX4308);
  and AND2_1514(WX4310,CRC_OUT_6_3,WX4883);
  and AND2_1515(WX4311,WX6380,WX4312);
  and AND2_1516(WX4314,WX4420,WX4883);
  and AND2_1517(WX4315,WX5087,WX4316);
  and AND2_1518(WX4320,WX4331,WX4882);
  and AND2_1519(WX4321,WX4327,WX4322);
  and AND2_1520(WX4324,CRC_OUT_6_2,WX4883);
  and AND2_1521(WX4325,WX6387,WX4326);
  and AND2_1522(WX4328,WX4422,WX4883);
  and AND2_1523(WX4329,WX5094,WX4330);
  and AND2_1524(WX4334,WX4345,WX4882);
  and AND2_1525(WX4335,WX4341,WX4336);
  and AND2_1526(WX4338,CRC_OUT_6_1,WX4883);
  and AND2_1527(WX4339,WX6394,WX4340);
  and AND2_1528(WX4342,WX4424,WX4883);
  and AND2_1529(WX4343,WX5101,WX4344);
  and AND2_1530(WX4348,WX4359,WX4882);
  and AND2_1531(WX4349,WX4355,WX4350);
  and AND2_1532(WX4352,CRC_OUT_6_0,WX4883);
  and AND2_1533(WX4353,WX6401,WX4354);
  and AND2_1534(WX4356,WX4426,WX4883);
  and AND2_1535(WX4357,WX5108,WX4358);
  and AND2_1536(WX4363,WX4366,RESET);
  and AND2_1537(WX4365,WX4368,RESET);
  and AND2_1538(WX4367,WX4370,RESET);
  and AND2_1539(WX4369,WX4372,RESET);
  and AND2_1540(WX4371,WX4374,RESET);
  and AND2_1541(WX4373,WX4376,RESET);
  and AND2_1542(WX4375,WX4378,RESET);
  and AND2_1543(WX4377,WX4380,RESET);
  and AND2_1544(WX4379,WX4382,RESET);
  and AND2_1545(WX4381,WX4384,RESET);
  and AND2_1546(WX4383,WX4386,RESET);
  and AND2_1547(WX4385,WX4388,RESET);
  and AND2_1548(WX4387,WX4390,RESET);
  and AND2_1549(WX4389,WX4392,RESET);
  and AND2_1550(WX4391,WX4394,RESET);
  and AND2_1551(WX4393,WX4396,RESET);
  and AND2_1552(WX4395,WX4398,RESET);
  and AND2_1553(WX4397,WX4400,RESET);
  and AND2_1554(WX4399,WX4402,RESET);
  and AND2_1555(WX4401,WX4404,RESET);
  and AND2_1556(WX4403,WX4406,RESET);
  and AND2_1557(WX4405,WX4408,RESET);
  and AND2_1558(WX4407,WX4410,RESET);
  and AND2_1559(WX4409,WX4412,RESET);
  and AND2_1560(WX4411,WX4414,RESET);
  and AND2_1561(WX4413,WX4416,RESET);
  and AND2_1562(WX4415,WX4418,RESET);
  and AND2_1563(WX4417,WX4420,RESET);
  and AND2_1564(WX4419,WX4422,RESET);
  and AND2_1565(WX4421,WX4424,RESET);
  and AND2_1566(WX4423,WX4426,RESET);
  and AND2_1567(WX4425,WX4362,RESET);
  and AND2_1568(WX4523,WX3927,RESET);
  and AND2_1569(WX4525,WX3941,RESET);
  and AND2_1570(WX4527,WX3955,RESET);
  and AND2_1571(WX4529,WX3969,RESET);
  and AND2_1572(WX4531,WX3983,RESET);
  and AND2_1573(WX4533,WX3997,RESET);
  and AND2_1574(WX4535,WX4011,RESET);
  and AND2_1575(WX4537,WX4025,RESET);
  and AND2_1576(WX4539,WX4039,RESET);
  and AND2_1577(WX4541,WX4053,RESET);
  and AND2_1578(WX4543,WX4067,RESET);
  and AND2_1579(WX4545,WX4081,RESET);
  and AND2_1580(WX4547,WX4095,RESET);
  and AND2_1581(WX4549,WX4109,RESET);
  and AND2_1582(WX4551,WX4123,RESET);
  and AND2_1583(WX4553,WX4137,RESET);
  and AND2_1584(WX4555,WX4151,RESET);
  and AND2_1585(WX4557,WX4165,RESET);
  and AND2_1586(WX4559,WX4179,RESET);
  and AND2_1587(WX4561,WX4193,RESET);
  and AND2_1588(WX4563,WX4207,RESET);
  and AND2_1589(WX4565,WX4221,RESET);
  and AND2_1590(WX4567,WX4235,RESET);
  and AND2_1591(WX4569,WX4249,RESET);
  and AND2_1592(WX4571,WX4263,RESET);
  and AND2_1593(WX4573,WX4277,RESET);
  and AND2_1594(WX4575,WX4291,RESET);
  and AND2_1595(WX4577,WX4305,RESET);
  and AND2_1596(WX4579,WX4319,RESET);
  and AND2_1597(WX4581,WX4333,RESET);
  and AND2_1598(WX4583,WX4347,RESET);
  and AND2_1599(WX4585,WX4361,RESET);
  and AND2_1600(WX4587,WX4524,RESET);
  and AND2_1601(WX4589,WX4526,RESET);
  and AND2_1602(WX4591,WX4528,RESET);
  and AND2_1603(WX4593,WX4530,RESET);
  and AND2_1604(WX4595,WX4532,RESET);
  and AND2_1605(WX4597,WX4534,RESET);
  and AND2_1606(WX4599,WX4536,RESET);
  and AND2_1607(WX4601,WX4538,RESET);
  and AND2_1608(WX4603,WX4540,RESET);
  and AND2_1609(WX4605,WX4542,RESET);
  and AND2_1610(WX4607,WX4544,RESET);
  and AND2_1611(WX4609,WX4546,RESET);
  and AND2_1612(WX4611,WX4548,RESET);
  and AND2_1613(WX4613,WX4550,RESET);
  and AND2_1614(WX4615,WX4552,RESET);
  and AND2_1615(WX4617,WX4554,RESET);
  and AND2_1616(WX4619,WX4556,RESET);
  and AND2_1617(WX4621,WX4558,RESET);
  and AND2_1618(WX4623,WX4560,RESET);
  and AND2_1619(WX4625,WX4562,RESET);
  and AND2_1620(WX4627,WX4564,RESET);
  and AND2_1621(WX4629,WX4566,RESET);
  and AND2_1622(WX4631,WX4568,RESET);
  and AND2_1623(WX4633,WX4570,RESET);
  and AND2_1624(WX4635,WX4572,RESET);
  and AND2_1625(WX4637,WX4574,RESET);
  and AND2_1626(WX4639,WX4576,RESET);
  and AND2_1627(WX4641,WX4578,RESET);
  and AND2_1628(WX4643,WX4580,RESET);
  and AND2_1629(WX4645,WX4582,RESET);
  and AND2_1630(WX4647,WX4584,RESET);
  and AND2_1631(WX4649,WX4586,RESET);
  and AND2_1632(WX4651,WX4588,RESET);
  and AND2_1633(WX4653,WX4590,RESET);
  and AND2_1634(WX4655,WX4592,RESET);
  and AND2_1635(WX4657,WX4594,RESET);
  and AND2_1636(WX4659,WX4596,RESET);
  and AND2_1637(WX4661,WX4598,RESET);
  and AND2_1638(WX4663,WX4600,RESET);
  and AND2_1639(WX4665,WX4602,RESET);
  and AND2_1640(WX4667,WX4604,RESET);
  and AND2_1641(WX4669,WX4606,RESET);
  and AND2_1642(WX4671,WX4608,RESET);
  and AND2_1643(WX4673,WX4610,RESET);
  and AND2_1644(WX4675,WX4612,RESET);
  and AND2_1645(WX4677,WX4614,RESET);
  and AND2_1646(WX4679,WX4616,RESET);
  and AND2_1647(WX4681,WX4618,RESET);
  and AND2_1648(WX4683,WX4620,RESET);
  and AND2_1649(WX4685,WX4622,RESET);
  and AND2_1650(WX4687,WX4624,RESET);
  and AND2_1651(WX4689,WX4626,RESET);
  and AND2_1652(WX4691,WX4628,RESET);
  and AND2_1653(WX4693,WX4630,RESET);
  and AND2_1654(WX4695,WX4632,RESET);
  and AND2_1655(WX4697,WX4634,RESET);
  and AND2_1656(WX4699,WX4636,RESET);
  and AND2_1657(WX4701,WX4638,RESET);
  and AND2_1658(WX4703,WX4640,RESET);
  and AND2_1659(WX4705,WX4642,RESET);
  and AND2_1660(WX4707,WX4644,RESET);
  and AND2_1661(WX4709,WX4646,RESET);
  and AND2_1662(WX4711,WX4648,RESET);
  and AND2_1663(WX4713,WX4650,RESET);
  and AND2_1664(WX4715,WX4652,RESET);
  and AND2_1665(WX4717,WX4654,RESET);
  and AND2_1666(WX4719,WX4656,RESET);
  and AND2_1667(WX4721,WX4658,RESET);
  and AND2_1668(WX4723,WX4660,RESET);
  and AND2_1669(WX4725,WX4662,RESET);
  and AND2_1670(WX4727,WX4664,RESET);
  and AND2_1671(WX4729,WX4666,RESET);
  and AND2_1672(WX4731,WX4668,RESET);
  and AND2_1673(WX4733,WX4670,RESET);
  and AND2_1674(WX4735,WX4672,RESET);
  and AND2_1675(WX4737,WX4674,RESET);
  and AND2_1676(WX4739,WX4676,RESET);
  and AND2_1677(WX4741,WX4678,RESET);
  and AND2_1678(WX4743,WX4680,RESET);
  and AND2_1679(WX4745,WX4682,RESET);
  and AND2_1680(WX4747,WX4684,RESET);
  and AND2_1681(WX4749,WX4686,RESET);
  and AND2_1682(WX4751,WX4688,RESET);
  and AND2_1683(WX4753,WX4690,RESET);
  and AND2_1684(WX4755,WX4692,RESET);
  and AND2_1685(WX4757,WX4694,RESET);
  and AND2_1686(WX4759,WX4696,RESET);
  and AND2_1687(WX4761,WX4698,RESET);
  and AND2_1688(WX4763,WX4700,RESET);
  and AND2_1689(WX4765,WX4702,RESET);
  and AND2_1690(WX4767,WX4704,RESET);
  and AND2_1691(WX4769,WX4706,RESET);
  and AND2_1692(WX4771,WX4708,RESET);
  and AND2_1693(WX4773,WX4710,RESET);
  and AND2_1694(WX4775,WX4712,RESET);
  and AND2_1695(WX4777,WX4714,RESET);
  and AND2_1696(WX4886,WX4885,WX4884);
  and AND2_1697(WX4887,WX4459,WX4888);
  and AND2_1698(WX4893,WX4892,WX4884);
  and AND2_1699(WX4894,WX4460,WX4895);
  and AND2_1700(WX4900,WX4899,WX4884);
  and AND2_1701(WX4901,WX4461,WX4902);
  and AND2_1702(WX4907,WX4906,WX4884);
  and AND2_1703(WX4908,WX4462,WX4909);
  and AND2_1704(WX4914,WX4913,WX4884);
  and AND2_1705(WX4915,WX4463,WX4916);
  and AND2_1706(WX4921,WX4920,WX4884);
  and AND2_1707(WX4922,WX4464,WX4923);
  and AND2_1708(WX4928,WX4927,WX4884);
  and AND2_1709(WX4929,WX4465,WX4930);
  and AND2_1710(WX4935,WX4934,WX4884);
  and AND2_1711(WX4936,WX4466,WX4937);
  and AND2_1712(WX4942,WX4941,WX4884);
  and AND2_1713(WX4943,WX4467,WX4944);
  and AND2_1714(WX4949,WX4948,WX4884);
  and AND2_1715(WX4950,WX4468,WX4951);
  and AND2_1716(WX4956,WX4955,WX4884);
  and AND2_1717(WX4957,WX4469,WX4958);
  and AND2_1718(WX4963,WX4962,WX4884);
  and AND2_1719(WX4964,WX4470,WX4965);
  and AND2_1720(WX4970,WX4969,WX4884);
  and AND2_1721(WX4971,WX4471,WX4972);
  and AND2_1722(WX4977,WX4976,WX4884);
  and AND2_1723(WX4978,WX4472,WX4979);
  and AND2_1724(WX4984,WX4983,WX4884);
  and AND2_1725(WX4985,WX4473,WX4986);
  and AND2_1726(WX4991,WX4990,WX4884);
  and AND2_1727(WX4992,WX4474,WX4993);
  and AND2_1728(WX4998,WX4997,WX4884);
  and AND2_1729(WX4999,WX4475,WX5000);
  and AND2_1730(WX5005,WX5004,WX4884);
  and AND2_1731(WX5006,WX4476,WX5007);
  and AND2_1732(WX5012,WX5011,WX4884);
  and AND2_1733(WX5013,WX4477,WX5014);
  and AND2_1734(WX5019,WX5018,WX4884);
  and AND2_1735(WX5020,WX4478,WX5021);
  and AND2_1736(WX5026,WX5025,WX4884);
  and AND2_1737(WX5027,WX4479,WX5028);
  and AND2_1738(WX5033,WX5032,WX4884);
  and AND2_1739(WX5034,WX4480,WX5035);
  and AND2_1740(WX5040,WX5039,WX4884);
  and AND2_1741(WX5041,WX4481,WX5042);
  and AND2_1742(WX5047,WX5046,WX4884);
  and AND2_1743(WX5048,WX4482,WX5049);
  and AND2_1744(WX5054,WX5053,WX4884);
  and AND2_1745(WX5055,WX4483,WX5056);
  and AND2_1746(WX5061,WX5060,WX4884);
  and AND2_1747(WX5062,WX4484,WX5063);
  and AND2_1748(WX5068,WX5067,WX4884);
  and AND2_1749(WX5069,WX4485,WX5070);
  and AND2_1750(WX5075,WX5074,WX4884);
  and AND2_1751(WX5076,WX4486,WX5077);
  and AND2_1752(WX5082,WX5081,WX4884);
  and AND2_1753(WX5083,WX4487,WX5084);
  and AND2_1754(WX5089,WX5088,WX4884);
  and AND2_1755(WX5090,WX4488,WX5091);
  and AND2_1756(WX5096,WX5095,WX4884);
  and AND2_1757(WX5097,WX4489,WX5098);
  and AND2_1758(WX5103,WX5102,WX4884);
  and AND2_1759(WX5104,WX4490,WX5105);
  and AND2_1760(WX5143,WX5113,WX5142);
  and AND2_1761(WX5145,WX5141,WX5142);
  and AND2_1762(WX5147,WX5140,WX5142);
  and AND2_1763(WX5149,WX5139,WX5142);
  and AND2_1764(WX5151,WX5112,WX5142);
  and AND2_1765(WX5153,WX5138,WX5142);
  and AND2_1766(WX5155,WX5137,WX5142);
  and AND2_1767(WX5157,WX5136,WX5142);
  and AND2_1768(WX5159,WX5135,WX5142);
  and AND2_1769(WX5161,WX5134,WX5142);
  and AND2_1770(WX5163,WX5133,WX5142);
  and AND2_1771(WX5165,WX5111,WX5142);
  and AND2_1772(WX5167,WX5132,WX5142);
  and AND2_1773(WX5169,WX5131,WX5142);
  and AND2_1774(WX5171,WX5130,WX5142);
  and AND2_1775(WX5173,WX5129,WX5142);
  and AND2_1776(WX5175,WX5110,WX5142);
  and AND2_1777(WX5177,WX5128,WX5142);
  and AND2_1778(WX5179,WX5127,WX5142);
  and AND2_1779(WX5181,WX5126,WX5142);
  and AND2_1780(WX5183,WX5125,WX5142);
  and AND2_1781(WX5185,WX5124,WX5142);
  and AND2_1782(WX5187,WX5123,WX5142);
  and AND2_1783(WX5189,WX5122,WX5142);
  and AND2_1784(WX5191,WX5121,WX5142);
  and AND2_1785(WX5193,WX5120,WX5142);
  and AND2_1786(WX5195,WX5119,WX5142);
  and AND2_1787(WX5197,WX5118,WX5142);
  and AND2_1788(WX5199,WX5117,WX5142);
  and AND2_1789(WX5201,WX5116,WX5142);
  and AND2_1790(WX5203,WX5115,WX5142);
  and AND2_1791(WX5205,WX5114,WX5142);
  and AND2_1792(WX5207,WX5218,WX6175);
  and AND2_1793(WX5208,WX5214,WX5209);
  and AND2_1794(WX5211,CRC_OUT_5_31,WX6176);
  and AND2_1795(WX5212,WX7477,WX5213);
  and AND2_1796(WX5215,WX5657,WX6176);
  and AND2_1797(WX5216,WX6184,WX5217);
  and AND2_1798(WX5221,WX5232,WX6175);
  and AND2_1799(WX5222,WX5228,WX5223);
  and AND2_1800(WX5225,CRC_OUT_5_30,WX6176);
  and AND2_1801(WX5226,WX7484,WX5227);
  and AND2_1802(WX5229,WX5659,WX6176);
  and AND2_1803(WX5230,WX6191,WX5231);
  and AND2_1804(WX5235,WX5246,WX6175);
  and AND2_1805(WX5236,WX5242,WX5237);
  and AND2_1806(WX5239,CRC_OUT_5_29,WX6176);
  and AND2_1807(WX5240,WX7491,WX5241);
  and AND2_1808(WX5243,WX5661,WX6176);
  and AND2_1809(WX5244,WX6198,WX5245);
  and AND2_1810(WX5249,WX5260,WX6175);
  and AND2_1811(WX5250,WX5256,WX5251);
  and AND2_1812(WX5253,CRC_OUT_5_28,WX6176);
  and AND2_1813(WX5254,WX7498,WX5255);
  and AND2_1814(WX5257,WX5663,WX6176);
  and AND2_1815(WX5258,WX6205,WX5259);
  and AND2_1816(WX5263,WX5274,WX6175);
  and AND2_1817(WX5264,WX5270,WX5265);
  and AND2_1818(WX5267,CRC_OUT_5_27,WX6176);
  and AND2_1819(WX5268,WX7505,WX5269);
  and AND2_1820(WX5271,WX5665,WX6176);
  and AND2_1821(WX5272,WX6212,WX5273);
  and AND2_1822(WX5277,WX5288,WX6175);
  and AND2_1823(WX5278,WX5284,WX5279);
  and AND2_1824(WX5281,CRC_OUT_5_26,WX6176);
  and AND2_1825(WX5282,WX7512,WX5283);
  and AND2_1826(WX5285,WX5667,WX6176);
  and AND2_1827(WX5286,WX6219,WX5287);
  and AND2_1828(WX5291,WX5302,WX6175);
  and AND2_1829(WX5292,WX5298,WX5293);
  and AND2_1830(WX5295,CRC_OUT_5_25,WX6176);
  and AND2_1831(WX5296,WX7519,WX5297);
  and AND2_1832(WX5299,WX5669,WX6176);
  and AND2_1833(WX5300,WX6226,WX5301);
  and AND2_1834(WX5305,WX5316,WX6175);
  and AND2_1835(WX5306,WX5312,WX5307);
  and AND2_1836(WX5309,CRC_OUT_5_24,WX6176);
  and AND2_1837(WX5310,WX7526,WX5311);
  and AND2_1838(WX5313,WX5671,WX6176);
  and AND2_1839(WX5314,WX6233,WX5315);
  and AND2_1840(WX5319,WX5330,WX6175);
  and AND2_1841(WX5320,WX5326,WX5321);
  and AND2_1842(WX5323,CRC_OUT_5_23,WX6176);
  and AND2_1843(WX5324,WX7533,WX5325);
  and AND2_1844(WX5327,WX5673,WX6176);
  and AND2_1845(WX5328,WX6240,WX5329);
  and AND2_1846(WX5333,WX5344,WX6175);
  and AND2_1847(WX5334,WX5340,WX5335);
  and AND2_1848(WX5337,CRC_OUT_5_22,WX6176);
  and AND2_1849(WX5338,WX7540,WX5339);
  and AND2_1850(WX5341,WX5675,WX6176);
  and AND2_1851(WX5342,WX6247,WX5343);
  and AND2_1852(WX5347,WX5358,WX6175);
  and AND2_1853(WX5348,WX5354,WX5349);
  and AND2_1854(WX5351,CRC_OUT_5_21,WX6176);
  and AND2_1855(WX5352,WX7547,WX5353);
  and AND2_1856(WX5355,WX5677,WX6176);
  and AND2_1857(WX5356,WX6254,WX5357);
  and AND2_1858(WX5361,WX5372,WX6175);
  and AND2_1859(WX5362,WX5368,WX5363);
  and AND2_1860(WX5365,CRC_OUT_5_20,WX6176);
  and AND2_1861(WX5366,WX7554,WX5367);
  and AND2_1862(WX5369,WX5679,WX6176);
  and AND2_1863(WX5370,WX6261,WX5371);
  and AND2_1864(WX5375,WX5386,WX6175);
  and AND2_1865(WX5376,WX5382,WX5377);
  and AND2_1866(WX5379,CRC_OUT_5_19,WX6176);
  and AND2_1867(WX5380,WX7561,WX5381);
  and AND2_1868(WX5383,WX5681,WX6176);
  and AND2_1869(WX5384,WX6268,WX5385);
  and AND2_1870(WX5389,WX5400,WX6175);
  and AND2_1871(WX5390,WX5396,WX5391);
  and AND2_1872(WX5393,CRC_OUT_5_18,WX6176);
  and AND2_1873(WX5394,WX7568,WX5395);
  and AND2_1874(WX5397,WX5683,WX6176);
  and AND2_1875(WX5398,WX6275,WX5399);
  and AND2_1876(WX5403,WX5414,WX6175);
  and AND2_1877(WX5404,WX5410,WX5405);
  and AND2_1878(WX5407,CRC_OUT_5_17,WX6176);
  and AND2_1879(WX5408,WX7575,WX5409);
  and AND2_1880(WX5411,WX5685,WX6176);
  and AND2_1881(WX5412,WX6282,WX5413);
  and AND2_1882(WX5417,WX5428,WX6175);
  and AND2_1883(WX5418,WX5424,WX5419);
  and AND2_1884(WX5421,CRC_OUT_5_16,WX6176);
  and AND2_1885(WX5422,WX7582,WX5423);
  and AND2_1886(WX5425,WX5687,WX6176);
  and AND2_1887(WX5426,WX6289,WX5427);
  and AND2_1888(WX5431,WX5442,WX6175);
  and AND2_1889(WX5432,WX5438,WX5433);
  and AND2_1890(WX5435,CRC_OUT_5_15,WX6176);
  and AND2_1891(WX5436,WX7589,WX5437);
  and AND2_1892(WX5439,WX5689,WX6176);
  and AND2_1893(WX5440,WX6296,WX5441);
  and AND2_1894(WX5445,WX5456,WX6175);
  and AND2_1895(WX5446,WX5452,WX5447);
  and AND2_1896(WX5449,CRC_OUT_5_14,WX6176);
  and AND2_1897(WX5450,WX7596,WX5451);
  and AND2_1898(WX5453,WX5691,WX6176);
  and AND2_1899(WX5454,WX6303,WX5455);
  and AND2_1900(WX5459,WX5470,WX6175);
  and AND2_1901(WX5460,WX5466,WX5461);
  and AND2_1902(WX5463,CRC_OUT_5_13,WX6176);
  and AND2_1903(WX5464,WX7603,WX5465);
  and AND2_1904(WX5467,WX5693,WX6176);
  and AND2_1905(WX5468,WX6310,WX5469);
  and AND2_1906(WX5473,WX5484,WX6175);
  and AND2_1907(WX5474,WX5480,WX5475);
  and AND2_1908(WX5477,CRC_OUT_5_12,WX6176);
  and AND2_1909(WX5478,WX7610,WX5479);
  and AND2_1910(WX5481,WX5695,WX6176);
  and AND2_1911(WX5482,WX6317,WX5483);
  and AND2_1912(WX5487,WX5498,WX6175);
  and AND2_1913(WX5488,WX5494,WX5489);
  and AND2_1914(WX5491,CRC_OUT_5_11,WX6176);
  and AND2_1915(WX5492,WX7617,WX5493);
  and AND2_1916(WX5495,WX5697,WX6176);
  and AND2_1917(WX5496,WX6324,WX5497);
  and AND2_1918(WX5501,WX5512,WX6175);
  and AND2_1919(WX5502,WX5508,WX5503);
  and AND2_1920(WX5505,CRC_OUT_5_10,WX6176);
  and AND2_1921(WX5506,WX7624,WX5507);
  and AND2_1922(WX5509,WX5699,WX6176);
  and AND2_1923(WX5510,WX6331,WX5511);
  and AND2_1924(WX5515,WX5526,WX6175);
  and AND2_1925(WX5516,WX5522,WX5517);
  and AND2_1926(WX5519,CRC_OUT_5_9,WX6176);
  and AND2_1927(WX5520,WX7631,WX5521);
  and AND2_1928(WX5523,WX5701,WX6176);
  and AND2_1929(WX5524,WX6338,WX5525);
  and AND2_1930(WX5529,WX5540,WX6175);
  and AND2_1931(WX5530,WX5536,WX5531);
  and AND2_1932(WX5533,CRC_OUT_5_8,WX6176);
  and AND2_1933(WX5534,WX7638,WX5535);
  and AND2_1934(WX5537,WX5703,WX6176);
  and AND2_1935(WX5538,WX6345,WX5539);
  and AND2_1936(WX5543,WX5554,WX6175);
  and AND2_1937(WX5544,WX5550,WX5545);
  and AND2_1938(WX5547,CRC_OUT_5_7,WX6176);
  and AND2_1939(WX5548,WX7645,WX5549);
  and AND2_1940(WX5551,WX5705,WX6176);
  and AND2_1941(WX5552,WX6352,WX5553);
  and AND2_1942(WX5557,WX5568,WX6175);
  and AND2_1943(WX5558,WX5564,WX5559);
  and AND2_1944(WX5561,CRC_OUT_5_6,WX6176);
  and AND2_1945(WX5562,WX7652,WX5563);
  and AND2_1946(WX5565,WX5707,WX6176);
  and AND2_1947(WX5566,WX6359,WX5567);
  and AND2_1948(WX5571,WX5582,WX6175);
  and AND2_1949(WX5572,WX5578,WX5573);
  and AND2_1950(WX5575,CRC_OUT_5_5,WX6176);
  and AND2_1951(WX5576,WX7659,WX5577);
  and AND2_1952(WX5579,WX5709,WX6176);
  and AND2_1953(WX5580,WX6366,WX5581);
  and AND2_1954(WX5585,WX5596,WX6175);
  and AND2_1955(WX5586,WX5592,WX5587);
  and AND2_1956(WX5589,CRC_OUT_5_4,WX6176);
  and AND2_1957(WX5590,WX7666,WX5591);
  and AND2_1958(WX5593,WX5711,WX6176);
  and AND2_1959(WX5594,WX6373,WX5595);
  and AND2_1960(WX5599,WX5610,WX6175);
  and AND2_1961(WX5600,WX5606,WX5601);
  and AND2_1962(WX5603,CRC_OUT_5_3,WX6176);
  and AND2_1963(WX5604,WX7673,WX5605);
  and AND2_1964(WX5607,WX5713,WX6176);
  and AND2_1965(WX5608,WX6380,WX5609);
  and AND2_1966(WX5613,WX5624,WX6175);
  and AND2_1967(WX5614,WX5620,WX5615);
  and AND2_1968(WX5617,CRC_OUT_5_2,WX6176);
  and AND2_1969(WX5618,WX7680,WX5619);
  and AND2_1970(WX5621,WX5715,WX6176);
  and AND2_1971(WX5622,WX6387,WX5623);
  and AND2_1972(WX5627,WX5638,WX6175);
  and AND2_1973(WX5628,WX5634,WX5629);
  and AND2_1974(WX5631,CRC_OUT_5_1,WX6176);
  and AND2_1975(WX5632,WX7687,WX5633);
  and AND2_1976(WX5635,WX5717,WX6176);
  and AND2_1977(WX5636,WX6394,WX5637);
  and AND2_1978(WX5641,WX5652,WX6175);
  and AND2_1979(WX5642,WX5648,WX5643);
  and AND2_1980(WX5645,CRC_OUT_5_0,WX6176);
  and AND2_1981(WX5646,WX7694,WX5647);
  and AND2_1982(WX5649,WX5719,WX6176);
  and AND2_1983(WX5650,WX6401,WX5651);
  and AND2_1984(WX5656,WX5659,RESET);
  and AND2_1985(WX5658,WX5661,RESET);
  and AND2_1986(WX5660,WX5663,RESET);
  and AND2_1987(WX5662,WX5665,RESET);
  and AND2_1988(WX5664,WX5667,RESET);
  and AND2_1989(WX5666,WX5669,RESET);
  and AND2_1990(WX5668,WX5671,RESET);
  and AND2_1991(WX5670,WX5673,RESET);
  and AND2_1992(WX5672,WX5675,RESET);
  and AND2_1993(WX5674,WX5677,RESET);
  and AND2_1994(WX5676,WX5679,RESET);
  and AND2_1995(WX5678,WX5681,RESET);
  and AND2_1996(WX5680,WX5683,RESET);
  and AND2_1997(WX5682,WX5685,RESET);
  and AND2_1998(WX5684,WX5687,RESET);
  and AND2_1999(WX5686,WX5689,RESET);
  and AND2_2000(WX5688,WX5691,RESET);
  and AND2_2001(WX5690,WX5693,RESET);
  and AND2_2002(WX5692,WX5695,RESET);
  and AND2_2003(WX5694,WX5697,RESET);
  and AND2_2004(WX5696,WX5699,RESET);
  and AND2_2005(WX5698,WX5701,RESET);
  and AND2_2006(WX5700,WX5703,RESET);
  and AND2_2007(WX5702,WX5705,RESET);
  and AND2_2008(WX5704,WX5707,RESET);
  and AND2_2009(WX5706,WX5709,RESET);
  and AND2_2010(WX5708,WX5711,RESET);
  and AND2_2011(WX5710,WX5713,RESET);
  and AND2_2012(WX5712,WX5715,RESET);
  and AND2_2013(WX5714,WX5717,RESET);
  and AND2_2014(WX5716,WX5719,RESET);
  and AND2_2015(WX5718,WX5655,RESET);
  and AND2_2016(WX5816,WX5220,RESET);
  and AND2_2017(WX5818,WX5234,RESET);
  and AND2_2018(WX5820,WX5248,RESET);
  and AND2_2019(WX5822,WX5262,RESET);
  and AND2_2020(WX5824,WX5276,RESET);
  and AND2_2021(WX5826,WX5290,RESET);
  and AND2_2022(WX5828,WX5304,RESET);
  and AND2_2023(WX5830,WX5318,RESET);
  and AND2_2024(WX5832,WX5332,RESET);
  and AND2_2025(WX5834,WX5346,RESET);
  and AND2_2026(WX5836,WX5360,RESET);
  and AND2_2027(WX5838,WX5374,RESET);
  and AND2_2028(WX5840,WX5388,RESET);
  and AND2_2029(WX5842,WX5402,RESET);
  and AND2_2030(WX5844,WX5416,RESET);
  and AND2_2031(WX5846,WX5430,RESET);
  and AND2_2032(WX5848,WX5444,RESET);
  and AND2_2033(WX5850,WX5458,RESET);
  and AND2_2034(WX5852,WX5472,RESET);
  and AND2_2035(WX5854,WX5486,RESET);
  and AND2_2036(WX5856,WX5500,RESET);
  and AND2_2037(WX5858,WX5514,RESET);
  and AND2_2038(WX5860,WX5528,RESET);
  and AND2_2039(WX5862,WX5542,RESET);
  and AND2_2040(WX5864,WX5556,RESET);
  and AND2_2041(WX5866,WX5570,RESET);
  and AND2_2042(WX5868,WX5584,RESET);
  and AND2_2043(WX5870,WX5598,RESET);
  and AND2_2044(WX5872,WX5612,RESET);
  and AND2_2045(WX5874,WX5626,RESET);
  and AND2_2046(WX5876,WX5640,RESET);
  and AND2_2047(WX5878,WX5654,RESET);
  and AND2_2048(WX5880,WX5817,RESET);
  and AND2_2049(WX5882,WX5819,RESET);
  and AND2_2050(WX5884,WX5821,RESET);
  and AND2_2051(WX5886,WX5823,RESET);
  and AND2_2052(WX5888,WX5825,RESET);
  and AND2_2053(WX5890,WX5827,RESET);
  and AND2_2054(WX5892,WX5829,RESET);
  and AND2_2055(WX5894,WX5831,RESET);
  and AND2_2056(WX5896,WX5833,RESET);
  and AND2_2057(WX5898,WX5835,RESET);
  and AND2_2058(WX5900,WX5837,RESET);
  and AND2_2059(WX5902,WX5839,RESET);
  and AND2_2060(WX5904,WX5841,RESET);
  and AND2_2061(WX5906,WX5843,RESET);
  and AND2_2062(WX5908,WX5845,RESET);
  and AND2_2063(WX5910,WX5847,RESET);
  and AND2_2064(WX5912,WX5849,RESET);
  and AND2_2065(WX5914,WX5851,RESET);
  and AND2_2066(WX5916,WX5853,RESET);
  and AND2_2067(WX5918,WX5855,RESET);
  and AND2_2068(WX5920,WX5857,RESET);
  and AND2_2069(WX5922,WX5859,RESET);
  and AND2_2070(WX5924,WX5861,RESET);
  and AND2_2071(WX5926,WX5863,RESET);
  and AND2_2072(WX5928,WX5865,RESET);
  and AND2_2073(WX5930,WX5867,RESET);
  and AND2_2074(WX5932,WX5869,RESET);
  and AND2_2075(WX5934,WX5871,RESET);
  and AND2_2076(WX5936,WX5873,RESET);
  and AND2_2077(WX5938,WX5875,RESET);
  and AND2_2078(WX5940,WX5877,RESET);
  and AND2_2079(WX5942,WX5879,RESET);
  and AND2_2080(WX5944,WX5881,RESET);
  and AND2_2081(WX5946,WX5883,RESET);
  and AND2_2082(WX5948,WX5885,RESET);
  and AND2_2083(WX5950,WX5887,RESET);
  and AND2_2084(WX5952,WX5889,RESET);
  and AND2_2085(WX5954,WX5891,RESET);
  and AND2_2086(WX5956,WX5893,RESET);
  and AND2_2087(WX5958,WX5895,RESET);
  and AND2_2088(WX5960,WX5897,RESET);
  and AND2_2089(WX5962,WX5899,RESET);
  and AND2_2090(WX5964,WX5901,RESET);
  and AND2_2091(WX5966,WX5903,RESET);
  and AND2_2092(WX5968,WX5905,RESET);
  and AND2_2093(WX5970,WX5907,RESET);
  and AND2_2094(WX5972,WX5909,RESET);
  and AND2_2095(WX5974,WX5911,RESET);
  and AND2_2096(WX5976,WX5913,RESET);
  and AND2_2097(WX5978,WX5915,RESET);
  and AND2_2098(WX5980,WX5917,RESET);
  and AND2_2099(WX5982,WX5919,RESET);
  and AND2_2100(WX5984,WX5921,RESET);
  and AND2_2101(WX5986,WX5923,RESET);
  and AND2_2102(WX5988,WX5925,RESET);
  and AND2_2103(WX5990,WX5927,RESET);
  and AND2_2104(WX5992,WX5929,RESET);
  and AND2_2105(WX5994,WX5931,RESET);
  and AND2_2106(WX5996,WX5933,RESET);
  and AND2_2107(WX5998,WX5935,RESET);
  and AND2_2108(WX6000,WX5937,RESET);
  and AND2_2109(WX6002,WX5939,RESET);
  and AND2_2110(WX6004,WX5941,RESET);
  and AND2_2111(WX6006,WX5943,RESET);
  and AND2_2112(WX6008,WX5945,RESET);
  and AND2_2113(WX6010,WX5947,RESET);
  and AND2_2114(WX6012,WX5949,RESET);
  and AND2_2115(WX6014,WX5951,RESET);
  and AND2_2116(WX6016,WX5953,RESET);
  and AND2_2117(WX6018,WX5955,RESET);
  and AND2_2118(WX6020,WX5957,RESET);
  and AND2_2119(WX6022,WX5959,RESET);
  and AND2_2120(WX6024,WX5961,RESET);
  and AND2_2121(WX6026,WX5963,RESET);
  and AND2_2122(WX6028,WX5965,RESET);
  and AND2_2123(WX6030,WX5967,RESET);
  and AND2_2124(WX6032,WX5969,RESET);
  and AND2_2125(WX6034,WX5971,RESET);
  and AND2_2126(WX6036,WX5973,RESET);
  and AND2_2127(WX6038,WX5975,RESET);
  and AND2_2128(WX6040,WX5977,RESET);
  and AND2_2129(WX6042,WX5979,RESET);
  and AND2_2130(WX6044,WX5981,RESET);
  and AND2_2131(WX6046,WX5983,RESET);
  and AND2_2132(WX6048,WX5985,RESET);
  and AND2_2133(WX6050,WX5987,RESET);
  and AND2_2134(WX6052,WX5989,RESET);
  and AND2_2135(WX6054,WX5991,RESET);
  and AND2_2136(WX6056,WX5993,RESET);
  and AND2_2137(WX6058,WX5995,RESET);
  and AND2_2138(WX6060,WX5997,RESET);
  and AND2_2139(WX6062,WX5999,RESET);
  and AND2_2140(WX6064,WX6001,RESET);
  and AND2_2141(WX6066,WX6003,RESET);
  and AND2_2142(WX6068,WX6005,RESET);
  and AND2_2143(WX6070,WX6007,RESET);
  and AND2_2144(WX6179,WX6178,WX6177);
  and AND2_2145(WX6180,WX5752,WX6181);
  and AND2_2146(WX6186,WX6185,WX6177);
  and AND2_2147(WX6187,WX5753,WX6188);
  and AND2_2148(WX6193,WX6192,WX6177);
  and AND2_2149(WX6194,WX5754,WX6195);
  and AND2_2150(WX6200,WX6199,WX6177);
  and AND2_2151(WX6201,WX5755,WX6202);
  and AND2_2152(WX6207,WX6206,WX6177);
  and AND2_2153(WX6208,WX5756,WX6209);
  and AND2_2154(WX6214,WX6213,WX6177);
  and AND2_2155(WX6215,WX5757,WX6216);
  and AND2_2156(WX6221,WX6220,WX6177);
  and AND2_2157(WX6222,WX5758,WX6223);
  and AND2_2158(WX6228,WX6227,WX6177);
  and AND2_2159(WX6229,WX5759,WX6230);
  and AND2_2160(WX6235,WX6234,WX6177);
  and AND2_2161(WX6236,WX5760,WX6237);
  and AND2_2162(WX6242,WX6241,WX6177);
  and AND2_2163(WX6243,WX5761,WX6244);
  and AND2_2164(WX6249,WX6248,WX6177);
  and AND2_2165(WX6250,WX5762,WX6251);
  and AND2_2166(WX6256,WX6255,WX6177);
  and AND2_2167(WX6257,WX5763,WX6258);
  and AND2_2168(WX6263,WX6262,WX6177);
  and AND2_2169(WX6264,WX5764,WX6265);
  and AND2_2170(WX6270,WX6269,WX6177);
  and AND2_2171(WX6271,WX5765,WX6272);
  and AND2_2172(WX6277,WX6276,WX6177);
  and AND2_2173(WX6278,WX5766,WX6279);
  and AND2_2174(WX6284,WX6283,WX6177);
  and AND2_2175(WX6285,WX5767,WX6286);
  and AND2_2176(WX6291,WX6290,WX6177);
  and AND2_2177(WX6292,WX5768,WX6293);
  and AND2_2178(WX6298,WX6297,WX6177);
  and AND2_2179(WX6299,WX5769,WX6300);
  and AND2_2180(WX6305,WX6304,WX6177);
  and AND2_2181(WX6306,WX5770,WX6307);
  and AND2_2182(WX6312,WX6311,WX6177);
  and AND2_2183(WX6313,WX5771,WX6314);
  and AND2_2184(WX6319,WX6318,WX6177);
  and AND2_2185(WX6320,WX5772,WX6321);
  and AND2_2186(WX6326,WX6325,WX6177);
  and AND2_2187(WX6327,WX5773,WX6328);
  and AND2_2188(WX6333,WX6332,WX6177);
  and AND2_2189(WX6334,WX5774,WX6335);
  and AND2_2190(WX6340,WX6339,WX6177);
  and AND2_2191(WX6341,WX5775,WX6342);
  and AND2_2192(WX6347,WX6346,WX6177);
  and AND2_2193(WX6348,WX5776,WX6349);
  and AND2_2194(WX6354,WX6353,WX6177);
  and AND2_2195(WX6355,WX5777,WX6356);
  and AND2_2196(WX6361,WX6360,WX6177);
  and AND2_2197(WX6362,WX5778,WX6363);
  and AND2_2198(WX6368,WX6367,WX6177);
  and AND2_2199(WX6369,WX5779,WX6370);
  and AND2_2200(WX6375,WX6374,WX6177);
  and AND2_2201(WX6376,WX5780,WX6377);
  and AND2_2202(WX6382,WX6381,WX6177);
  and AND2_2203(WX6383,WX5781,WX6384);
  and AND2_2204(WX6389,WX6388,WX6177);
  and AND2_2205(WX6390,WX5782,WX6391);
  and AND2_2206(WX6396,WX6395,WX6177);
  and AND2_2207(WX6397,WX5783,WX6398);
  and AND2_2208(WX6436,WX6406,WX6435);
  and AND2_2209(WX6438,WX6434,WX6435);
  and AND2_2210(WX6440,WX6433,WX6435);
  and AND2_2211(WX6442,WX6432,WX6435);
  and AND2_2212(WX6444,WX6405,WX6435);
  and AND2_2213(WX6446,WX6431,WX6435);
  and AND2_2214(WX6448,WX6430,WX6435);
  and AND2_2215(WX6450,WX6429,WX6435);
  and AND2_2216(WX6452,WX6428,WX6435);
  and AND2_2217(WX6454,WX6427,WX6435);
  and AND2_2218(WX6456,WX6426,WX6435);
  and AND2_2219(WX6458,WX6404,WX6435);
  and AND2_2220(WX6460,WX6425,WX6435);
  and AND2_2221(WX6462,WX6424,WX6435);
  and AND2_2222(WX6464,WX6423,WX6435);
  and AND2_2223(WX6466,WX6422,WX6435);
  and AND2_2224(WX6468,WX6403,WX6435);
  and AND2_2225(WX6470,WX6421,WX6435);
  and AND2_2226(WX6472,WX6420,WX6435);
  and AND2_2227(WX6474,WX6419,WX6435);
  and AND2_2228(WX6476,WX6418,WX6435);
  and AND2_2229(WX6478,WX6417,WX6435);
  and AND2_2230(WX6480,WX6416,WX6435);
  and AND2_2231(WX6482,WX6415,WX6435);
  and AND2_2232(WX6484,WX6414,WX6435);
  and AND2_2233(WX6486,WX6413,WX6435);
  and AND2_2234(WX6488,WX6412,WX6435);
  and AND2_2235(WX6490,WX6411,WX6435);
  and AND2_2236(WX6492,WX6410,WX6435);
  and AND2_2237(WX6494,WX6409,WX6435);
  and AND2_2238(WX6496,WX6408,WX6435);
  and AND2_2239(WX6498,WX6407,WX6435);
  and AND2_2240(WX6500,WX6511,WX7468);
  and AND2_2241(WX6501,WX6507,WX6502);
  and AND2_2242(WX6504,CRC_OUT_4_31,WX7469);
  and AND2_2243(WX6505,WX8770,WX6506);
  and AND2_2244(WX6508,WX6950,WX7469);
  and AND2_2245(WX6509,WX7477,WX6510);
  and AND2_2246(WX6514,WX6525,WX7468);
  and AND2_2247(WX6515,WX6521,WX6516);
  and AND2_2248(WX6518,CRC_OUT_4_30,WX7469);
  and AND2_2249(WX6519,WX8777,WX6520);
  and AND2_2250(WX6522,WX6952,WX7469);
  and AND2_2251(WX6523,WX7484,WX6524);
  and AND2_2252(WX6528,WX6539,WX7468);
  and AND2_2253(WX6529,WX6535,WX6530);
  and AND2_2254(WX6532,CRC_OUT_4_29,WX7469);
  and AND2_2255(WX6533,WX8784,WX6534);
  and AND2_2256(WX6536,WX6954,WX7469);
  and AND2_2257(WX6537,WX7491,WX6538);
  and AND2_2258(WX6542,WX6553,WX7468);
  and AND2_2259(WX6543,WX6549,WX6544);
  and AND2_2260(WX6546,CRC_OUT_4_28,WX7469);
  and AND2_2261(WX6547,WX8791,WX6548);
  and AND2_2262(WX6550,WX6956,WX7469);
  and AND2_2263(WX6551,WX7498,WX6552);
  and AND2_2264(WX6556,WX6567,WX7468);
  and AND2_2265(WX6557,WX6563,WX6558);
  and AND2_2266(WX6560,CRC_OUT_4_27,WX7469);
  and AND2_2267(WX6561,WX8798,WX6562);
  and AND2_2268(WX6564,WX6958,WX7469);
  and AND2_2269(WX6565,WX7505,WX6566);
  and AND2_2270(WX6570,WX6581,WX7468);
  and AND2_2271(WX6571,WX6577,WX6572);
  and AND2_2272(WX6574,CRC_OUT_4_26,WX7469);
  and AND2_2273(WX6575,WX8805,WX6576);
  and AND2_2274(WX6578,WX6960,WX7469);
  and AND2_2275(WX6579,WX7512,WX6580);
  and AND2_2276(WX6584,WX6595,WX7468);
  and AND2_2277(WX6585,WX6591,WX6586);
  and AND2_2278(WX6588,CRC_OUT_4_25,WX7469);
  and AND2_2279(WX6589,WX8812,WX6590);
  and AND2_2280(WX6592,WX6962,WX7469);
  and AND2_2281(WX6593,WX7519,WX6594);
  and AND2_2282(WX6598,WX6609,WX7468);
  and AND2_2283(WX6599,WX6605,WX6600);
  and AND2_2284(WX6602,CRC_OUT_4_24,WX7469);
  and AND2_2285(WX6603,WX8819,WX6604);
  and AND2_2286(WX6606,WX6964,WX7469);
  and AND2_2287(WX6607,WX7526,WX6608);
  and AND2_2288(WX6612,WX6623,WX7468);
  and AND2_2289(WX6613,WX6619,WX6614);
  and AND2_2290(WX6616,CRC_OUT_4_23,WX7469);
  and AND2_2291(WX6617,WX8826,WX6618);
  and AND2_2292(WX6620,WX6966,WX7469);
  and AND2_2293(WX6621,WX7533,WX6622);
  and AND2_2294(WX6626,WX6637,WX7468);
  and AND2_2295(WX6627,WX6633,WX6628);
  and AND2_2296(WX6630,CRC_OUT_4_22,WX7469);
  and AND2_2297(WX6631,WX8833,WX6632);
  and AND2_2298(WX6634,WX6968,WX7469);
  and AND2_2299(WX6635,WX7540,WX6636);
  and AND2_2300(WX6640,WX6651,WX7468);
  and AND2_2301(WX6641,WX6647,WX6642);
  and AND2_2302(WX6644,CRC_OUT_4_21,WX7469);
  and AND2_2303(WX6645,WX8840,WX6646);
  and AND2_2304(WX6648,WX6970,WX7469);
  and AND2_2305(WX6649,WX7547,WX6650);
  and AND2_2306(WX6654,WX6665,WX7468);
  and AND2_2307(WX6655,WX6661,WX6656);
  and AND2_2308(WX6658,CRC_OUT_4_20,WX7469);
  and AND2_2309(WX6659,WX8847,WX6660);
  and AND2_2310(WX6662,WX6972,WX7469);
  and AND2_2311(WX6663,WX7554,WX6664);
  and AND2_2312(WX6668,WX6679,WX7468);
  and AND2_2313(WX6669,WX6675,WX6670);
  and AND2_2314(WX6672,CRC_OUT_4_19,WX7469);
  and AND2_2315(WX6673,WX8854,WX6674);
  and AND2_2316(WX6676,WX6974,WX7469);
  and AND2_2317(WX6677,WX7561,WX6678);
  and AND2_2318(WX6682,WX6693,WX7468);
  and AND2_2319(WX6683,WX6689,WX6684);
  and AND2_2320(WX6686,CRC_OUT_4_18,WX7469);
  and AND2_2321(WX6687,WX8861,WX6688);
  and AND2_2322(WX6690,WX6976,WX7469);
  and AND2_2323(WX6691,WX7568,WX6692);
  and AND2_2324(WX6696,WX6707,WX7468);
  and AND2_2325(WX6697,WX6703,WX6698);
  and AND2_2326(WX6700,CRC_OUT_4_17,WX7469);
  and AND2_2327(WX6701,WX8868,WX6702);
  and AND2_2328(WX6704,WX6978,WX7469);
  and AND2_2329(WX6705,WX7575,WX6706);
  and AND2_2330(WX6710,WX6721,WX7468);
  and AND2_2331(WX6711,WX6717,WX6712);
  and AND2_2332(WX6714,CRC_OUT_4_16,WX7469);
  and AND2_2333(WX6715,WX8875,WX6716);
  and AND2_2334(WX6718,WX6980,WX7469);
  and AND2_2335(WX6719,WX7582,WX6720);
  and AND2_2336(WX6724,WX6735,WX7468);
  and AND2_2337(WX6725,WX6731,WX6726);
  and AND2_2338(WX6728,CRC_OUT_4_15,WX7469);
  and AND2_2339(WX6729,WX8882,WX6730);
  and AND2_2340(WX6732,WX6982,WX7469);
  and AND2_2341(WX6733,WX7589,WX6734);
  and AND2_2342(WX6738,WX6749,WX7468);
  and AND2_2343(WX6739,WX6745,WX6740);
  and AND2_2344(WX6742,CRC_OUT_4_14,WX7469);
  and AND2_2345(WX6743,WX8889,WX6744);
  and AND2_2346(WX6746,WX6984,WX7469);
  and AND2_2347(WX6747,WX7596,WX6748);
  and AND2_2348(WX6752,WX6763,WX7468);
  and AND2_2349(WX6753,WX6759,WX6754);
  and AND2_2350(WX6756,CRC_OUT_4_13,WX7469);
  and AND2_2351(WX6757,WX8896,WX6758);
  and AND2_2352(WX6760,WX6986,WX7469);
  and AND2_2353(WX6761,WX7603,WX6762);
  and AND2_2354(WX6766,WX6777,WX7468);
  and AND2_2355(WX6767,WX6773,WX6768);
  and AND2_2356(WX6770,CRC_OUT_4_12,WX7469);
  and AND2_2357(WX6771,WX8903,WX6772);
  and AND2_2358(WX6774,WX6988,WX7469);
  and AND2_2359(WX6775,WX7610,WX6776);
  and AND2_2360(WX6780,WX6791,WX7468);
  and AND2_2361(WX6781,WX6787,WX6782);
  and AND2_2362(WX6784,CRC_OUT_4_11,WX7469);
  and AND2_2363(WX6785,WX8910,WX6786);
  and AND2_2364(WX6788,WX6990,WX7469);
  and AND2_2365(WX6789,WX7617,WX6790);
  and AND2_2366(WX6794,WX6805,WX7468);
  and AND2_2367(WX6795,WX6801,WX6796);
  and AND2_2368(WX6798,CRC_OUT_4_10,WX7469);
  and AND2_2369(WX6799,WX8917,WX6800);
  and AND2_2370(WX6802,WX6992,WX7469);
  and AND2_2371(WX6803,WX7624,WX6804);
  and AND2_2372(WX6808,WX6819,WX7468);
  and AND2_2373(WX6809,WX6815,WX6810);
  and AND2_2374(WX6812,CRC_OUT_4_9,WX7469);
  and AND2_2375(WX6813,WX8924,WX6814);
  and AND2_2376(WX6816,WX6994,WX7469);
  and AND2_2377(WX6817,WX7631,WX6818);
  and AND2_2378(WX6822,WX6833,WX7468);
  and AND2_2379(WX6823,WX6829,WX6824);
  and AND2_2380(WX6826,CRC_OUT_4_8,WX7469);
  and AND2_2381(WX6827,WX8931,WX6828);
  and AND2_2382(WX6830,WX6996,WX7469);
  and AND2_2383(WX6831,WX7638,WX6832);
  and AND2_2384(WX6836,WX6847,WX7468);
  and AND2_2385(WX6837,WX6843,WX6838);
  and AND2_2386(WX6840,CRC_OUT_4_7,WX7469);
  and AND2_2387(WX6841,WX8938,WX6842);
  and AND2_2388(WX6844,WX6998,WX7469);
  and AND2_2389(WX6845,WX7645,WX6846);
  and AND2_2390(WX6850,WX6861,WX7468);
  and AND2_2391(WX6851,WX6857,WX6852);
  and AND2_2392(WX6854,CRC_OUT_4_6,WX7469);
  and AND2_2393(WX6855,WX8945,WX6856);
  and AND2_2394(WX6858,WX7000,WX7469);
  and AND2_2395(WX6859,WX7652,WX6860);
  and AND2_2396(WX6864,WX6875,WX7468);
  and AND2_2397(WX6865,WX6871,WX6866);
  and AND2_2398(WX6868,CRC_OUT_4_5,WX7469);
  and AND2_2399(WX6869,WX8952,WX6870);
  and AND2_2400(WX6872,WX7002,WX7469);
  and AND2_2401(WX6873,WX7659,WX6874);
  and AND2_2402(WX6878,WX6889,WX7468);
  and AND2_2403(WX6879,WX6885,WX6880);
  and AND2_2404(WX6882,CRC_OUT_4_4,WX7469);
  and AND2_2405(WX6883,WX8959,WX6884);
  and AND2_2406(WX6886,WX7004,WX7469);
  and AND2_2407(WX6887,WX7666,WX6888);
  and AND2_2408(WX6892,WX6903,WX7468);
  and AND2_2409(WX6893,WX6899,WX6894);
  and AND2_2410(WX6896,CRC_OUT_4_3,WX7469);
  and AND2_2411(WX6897,WX8966,WX6898);
  and AND2_2412(WX6900,WX7006,WX7469);
  and AND2_2413(WX6901,WX7673,WX6902);
  and AND2_2414(WX6906,WX6917,WX7468);
  and AND2_2415(WX6907,WX6913,WX6908);
  and AND2_2416(WX6910,CRC_OUT_4_2,WX7469);
  and AND2_2417(WX6911,WX8973,WX6912);
  and AND2_2418(WX6914,WX7008,WX7469);
  and AND2_2419(WX6915,WX7680,WX6916);
  and AND2_2420(WX6920,WX6931,WX7468);
  and AND2_2421(WX6921,WX6927,WX6922);
  and AND2_2422(WX6924,CRC_OUT_4_1,WX7469);
  and AND2_2423(WX6925,WX8980,WX6926);
  and AND2_2424(WX6928,WX7010,WX7469);
  and AND2_2425(WX6929,WX7687,WX6930);
  and AND2_2426(WX6934,WX6945,WX7468);
  and AND2_2427(WX6935,WX6941,WX6936);
  and AND2_2428(WX6938,CRC_OUT_4_0,WX7469);
  and AND2_2429(WX6939,WX8987,WX6940);
  and AND2_2430(WX6942,WX7012,WX7469);
  and AND2_2431(WX6943,WX7694,WX6944);
  and AND2_2432(WX6949,WX6952,RESET);
  and AND2_2433(WX6951,WX6954,RESET);
  and AND2_2434(WX6953,WX6956,RESET);
  and AND2_2435(WX6955,WX6958,RESET);
  and AND2_2436(WX6957,WX6960,RESET);
  and AND2_2437(WX6959,WX6962,RESET);
  and AND2_2438(WX6961,WX6964,RESET);
  and AND2_2439(WX6963,WX6966,RESET);
  and AND2_2440(WX6965,WX6968,RESET);
  and AND2_2441(WX6967,WX6970,RESET);
  and AND2_2442(WX6969,WX6972,RESET);
  and AND2_2443(WX6971,WX6974,RESET);
  and AND2_2444(WX6973,WX6976,RESET);
  and AND2_2445(WX6975,WX6978,RESET);
  and AND2_2446(WX6977,WX6980,RESET);
  and AND2_2447(WX6979,WX6982,RESET);
  and AND2_2448(WX6981,WX6984,RESET);
  and AND2_2449(WX6983,WX6986,RESET);
  and AND2_2450(WX6985,WX6988,RESET);
  and AND2_2451(WX6987,WX6990,RESET);
  and AND2_2452(WX6989,WX6992,RESET);
  and AND2_2453(WX6991,WX6994,RESET);
  and AND2_2454(WX6993,WX6996,RESET);
  and AND2_2455(WX6995,WX6998,RESET);
  and AND2_2456(WX6997,WX7000,RESET);
  and AND2_2457(WX6999,WX7002,RESET);
  and AND2_2458(WX7001,WX7004,RESET);
  and AND2_2459(WX7003,WX7006,RESET);
  and AND2_2460(WX7005,WX7008,RESET);
  and AND2_2461(WX7007,WX7010,RESET);
  and AND2_2462(WX7009,WX7012,RESET);
  and AND2_2463(WX7011,WX6948,RESET);
  and AND2_2464(WX7109,WX6513,RESET);
  and AND2_2465(WX7111,WX6527,RESET);
  and AND2_2466(WX7113,WX6541,RESET);
  and AND2_2467(WX7115,WX6555,RESET);
  and AND2_2468(WX7117,WX6569,RESET);
  and AND2_2469(WX7119,WX6583,RESET);
  and AND2_2470(WX7121,WX6597,RESET);
  and AND2_2471(WX7123,WX6611,RESET);
  and AND2_2472(WX7125,WX6625,RESET);
  and AND2_2473(WX7127,WX6639,RESET);
  and AND2_2474(WX7129,WX6653,RESET);
  and AND2_2475(WX7131,WX6667,RESET);
  and AND2_2476(WX7133,WX6681,RESET);
  and AND2_2477(WX7135,WX6695,RESET);
  and AND2_2478(WX7137,WX6709,RESET);
  and AND2_2479(WX7139,WX6723,RESET);
  and AND2_2480(WX7141,WX6737,RESET);
  and AND2_2481(WX7143,WX6751,RESET);
  and AND2_2482(WX7145,WX6765,RESET);
  and AND2_2483(WX7147,WX6779,RESET);
  and AND2_2484(WX7149,WX6793,RESET);
  and AND2_2485(WX7151,WX6807,RESET);
  and AND2_2486(WX7153,WX6821,RESET);
  and AND2_2487(WX7155,WX6835,RESET);
  and AND2_2488(WX7157,WX6849,RESET);
  and AND2_2489(WX7159,WX6863,RESET);
  and AND2_2490(WX7161,WX6877,RESET);
  and AND2_2491(WX7163,WX6891,RESET);
  and AND2_2492(WX7165,WX6905,RESET);
  and AND2_2493(WX7167,WX6919,RESET);
  and AND2_2494(WX7169,WX6933,RESET);
  and AND2_2495(WX7171,WX6947,RESET);
  and AND2_2496(WX7173,WX7110,RESET);
  and AND2_2497(WX7175,WX7112,RESET);
  and AND2_2498(WX7177,WX7114,RESET);
  and AND2_2499(WX7179,WX7116,RESET);
  and AND2_2500(WX7181,WX7118,RESET);
  and AND2_2501(WX7183,WX7120,RESET);
  and AND2_2502(WX7185,WX7122,RESET);
  and AND2_2503(WX7187,WX7124,RESET);
  and AND2_2504(WX7189,WX7126,RESET);
  and AND2_2505(WX7191,WX7128,RESET);
  and AND2_2506(WX7193,WX7130,RESET);
  and AND2_2507(WX7195,WX7132,RESET);
  and AND2_2508(WX7197,WX7134,RESET);
  and AND2_2509(WX7199,WX7136,RESET);
  and AND2_2510(WX7201,WX7138,RESET);
  and AND2_2511(WX7203,WX7140,RESET);
  and AND2_2512(WX7205,WX7142,RESET);
  and AND2_2513(WX7207,WX7144,RESET);
  and AND2_2514(WX7209,WX7146,RESET);
  and AND2_2515(WX7211,WX7148,RESET);
  and AND2_2516(WX7213,WX7150,RESET);
  and AND2_2517(WX7215,WX7152,RESET);
  and AND2_2518(WX7217,WX7154,RESET);
  and AND2_2519(WX7219,WX7156,RESET);
  and AND2_2520(WX7221,WX7158,RESET);
  and AND2_2521(WX7223,WX7160,RESET);
  and AND2_2522(WX7225,WX7162,RESET);
  and AND2_2523(WX7227,WX7164,RESET);
  and AND2_2524(WX7229,WX7166,RESET);
  and AND2_2525(WX7231,WX7168,RESET);
  and AND2_2526(WX7233,WX7170,RESET);
  and AND2_2527(WX7235,WX7172,RESET);
  and AND2_2528(WX7237,WX7174,RESET);
  and AND2_2529(WX7239,WX7176,RESET);
  and AND2_2530(WX7241,WX7178,RESET);
  and AND2_2531(WX7243,WX7180,RESET);
  and AND2_2532(WX7245,WX7182,RESET);
  and AND2_2533(WX7247,WX7184,RESET);
  and AND2_2534(WX7249,WX7186,RESET);
  and AND2_2535(WX7251,WX7188,RESET);
  and AND2_2536(WX7253,WX7190,RESET);
  and AND2_2537(WX7255,WX7192,RESET);
  and AND2_2538(WX7257,WX7194,RESET);
  and AND2_2539(WX7259,WX7196,RESET);
  and AND2_2540(WX7261,WX7198,RESET);
  and AND2_2541(WX7263,WX7200,RESET);
  and AND2_2542(WX7265,WX7202,RESET);
  and AND2_2543(WX7267,WX7204,RESET);
  and AND2_2544(WX7269,WX7206,RESET);
  and AND2_2545(WX7271,WX7208,RESET);
  and AND2_2546(WX7273,WX7210,RESET);
  and AND2_2547(WX7275,WX7212,RESET);
  and AND2_2548(WX7277,WX7214,RESET);
  and AND2_2549(WX7279,WX7216,RESET);
  and AND2_2550(WX7281,WX7218,RESET);
  and AND2_2551(WX7283,WX7220,RESET);
  and AND2_2552(WX7285,WX7222,RESET);
  and AND2_2553(WX7287,WX7224,RESET);
  and AND2_2554(WX7289,WX7226,RESET);
  and AND2_2555(WX7291,WX7228,RESET);
  and AND2_2556(WX7293,WX7230,RESET);
  and AND2_2557(WX7295,WX7232,RESET);
  and AND2_2558(WX7297,WX7234,RESET);
  and AND2_2559(WX7299,WX7236,RESET);
  and AND2_2560(WX7301,WX7238,RESET);
  and AND2_2561(WX7303,WX7240,RESET);
  and AND2_2562(WX7305,WX7242,RESET);
  and AND2_2563(WX7307,WX7244,RESET);
  and AND2_2564(WX7309,WX7246,RESET);
  and AND2_2565(WX7311,WX7248,RESET);
  and AND2_2566(WX7313,WX7250,RESET);
  and AND2_2567(WX7315,WX7252,RESET);
  and AND2_2568(WX7317,WX7254,RESET);
  and AND2_2569(WX7319,WX7256,RESET);
  and AND2_2570(WX7321,WX7258,RESET);
  and AND2_2571(WX7323,WX7260,RESET);
  and AND2_2572(WX7325,WX7262,RESET);
  and AND2_2573(WX7327,WX7264,RESET);
  and AND2_2574(WX7329,WX7266,RESET);
  and AND2_2575(WX7331,WX7268,RESET);
  and AND2_2576(WX7333,WX7270,RESET);
  and AND2_2577(WX7335,WX7272,RESET);
  and AND2_2578(WX7337,WX7274,RESET);
  and AND2_2579(WX7339,WX7276,RESET);
  and AND2_2580(WX7341,WX7278,RESET);
  and AND2_2581(WX7343,WX7280,RESET);
  and AND2_2582(WX7345,WX7282,RESET);
  and AND2_2583(WX7347,WX7284,RESET);
  and AND2_2584(WX7349,WX7286,RESET);
  and AND2_2585(WX7351,WX7288,RESET);
  and AND2_2586(WX7353,WX7290,RESET);
  and AND2_2587(WX7355,WX7292,RESET);
  and AND2_2588(WX7357,WX7294,RESET);
  and AND2_2589(WX7359,WX7296,RESET);
  and AND2_2590(WX7361,WX7298,RESET);
  and AND2_2591(WX7363,WX7300,RESET);
  and AND2_2592(WX7472,WX7471,WX7470);
  and AND2_2593(WX7473,WX7045,WX7474);
  and AND2_2594(WX7479,WX7478,WX7470);
  and AND2_2595(WX7480,WX7046,WX7481);
  and AND2_2596(WX7486,WX7485,WX7470);
  and AND2_2597(WX7487,WX7047,WX7488);
  and AND2_2598(WX7493,WX7492,WX7470);
  and AND2_2599(WX7494,WX7048,WX7495);
  and AND2_2600(WX7500,WX7499,WX7470);
  and AND2_2601(WX7501,WX7049,WX7502);
  and AND2_2602(WX7507,WX7506,WX7470);
  and AND2_2603(WX7508,WX7050,WX7509);
  and AND2_2604(WX7514,WX7513,WX7470);
  and AND2_2605(WX7515,WX7051,WX7516);
  and AND2_2606(WX7521,WX7520,WX7470);
  and AND2_2607(WX7522,WX7052,WX7523);
  and AND2_2608(WX7528,WX7527,WX7470);
  and AND2_2609(WX7529,WX7053,WX7530);
  and AND2_2610(WX7535,WX7534,WX7470);
  and AND2_2611(WX7536,WX7054,WX7537);
  and AND2_2612(WX7542,WX7541,WX7470);
  and AND2_2613(WX7543,WX7055,WX7544);
  and AND2_2614(WX7549,WX7548,WX7470);
  and AND2_2615(WX7550,WX7056,WX7551);
  and AND2_2616(WX7556,WX7555,WX7470);
  and AND2_2617(WX7557,WX7057,WX7558);
  and AND2_2618(WX7563,WX7562,WX7470);
  and AND2_2619(WX7564,WX7058,WX7565);
  and AND2_2620(WX7570,WX7569,WX7470);
  and AND2_2621(WX7571,WX7059,WX7572);
  and AND2_2622(WX7577,WX7576,WX7470);
  and AND2_2623(WX7578,WX7060,WX7579);
  and AND2_2624(WX7584,WX7583,WX7470);
  and AND2_2625(WX7585,WX7061,WX7586);
  and AND2_2626(WX7591,WX7590,WX7470);
  and AND2_2627(WX7592,WX7062,WX7593);
  and AND2_2628(WX7598,WX7597,WX7470);
  and AND2_2629(WX7599,WX7063,WX7600);
  and AND2_2630(WX7605,WX7604,WX7470);
  and AND2_2631(WX7606,WX7064,WX7607);
  and AND2_2632(WX7612,WX7611,WX7470);
  and AND2_2633(WX7613,WX7065,WX7614);
  and AND2_2634(WX7619,WX7618,WX7470);
  and AND2_2635(WX7620,WX7066,WX7621);
  and AND2_2636(WX7626,WX7625,WX7470);
  and AND2_2637(WX7627,WX7067,WX7628);
  and AND2_2638(WX7633,WX7632,WX7470);
  and AND2_2639(WX7634,WX7068,WX7635);
  and AND2_2640(WX7640,WX7639,WX7470);
  and AND2_2641(WX7641,WX7069,WX7642);
  and AND2_2642(WX7647,WX7646,WX7470);
  and AND2_2643(WX7648,WX7070,WX7649);
  and AND2_2644(WX7654,WX7653,WX7470);
  and AND2_2645(WX7655,WX7071,WX7656);
  and AND2_2646(WX7661,WX7660,WX7470);
  and AND2_2647(WX7662,WX7072,WX7663);
  and AND2_2648(WX7668,WX7667,WX7470);
  and AND2_2649(WX7669,WX7073,WX7670);
  and AND2_2650(WX7675,WX7674,WX7470);
  and AND2_2651(WX7676,WX7074,WX7677);
  and AND2_2652(WX7682,WX7681,WX7470);
  and AND2_2653(WX7683,WX7075,WX7684);
  and AND2_2654(WX7689,WX7688,WX7470);
  and AND2_2655(WX7690,WX7076,WX7691);
  and AND2_2656(WX7729,WX7699,WX7728);
  and AND2_2657(WX7731,WX7727,WX7728);
  and AND2_2658(WX7733,WX7726,WX7728);
  and AND2_2659(WX7735,WX7725,WX7728);
  and AND2_2660(WX7737,WX7698,WX7728);
  and AND2_2661(WX7739,WX7724,WX7728);
  and AND2_2662(WX7741,WX7723,WX7728);
  and AND2_2663(WX7743,WX7722,WX7728);
  and AND2_2664(WX7745,WX7721,WX7728);
  and AND2_2665(WX7747,WX7720,WX7728);
  and AND2_2666(WX7749,WX7719,WX7728);
  and AND2_2667(WX7751,WX7697,WX7728);
  and AND2_2668(WX7753,WX7718,WX7728);
  and AND2_2669(WX7755,WX7717,WX7728);
  and AND2_2670(WX7757,WX7716,WX7728);
  and AND2_2671(WX7759,WX7715,WX7728);
  and AND2_2672(WX7761,WX7696,WX7728);
  and AND2_2673(WX7763,WX7714,WX7728);
  and AND2_2674(WX7765,WX7713,WX7728);
  and AND2_2675(WX7767,WX7712,WX7728);
  and AND2_2676(WX7769,WX7711,WX7728);
  and AND2_2677(WX7771,WX7710,WX7728);
  and AND2_2678(WX7773,WX7709,WX7728);
  and AND2_2679(WX7775,WX7708,WX7728);
  and AND2_2680(WX7777,WX7707,WX7728);
  and AND2_2681(WX7779,WX7706,WX7728);
  and AND2_2682(WX7781,WX7705,WX7728);
  and AND2_2683(WX7783,WX7704,WX7728);
  and AND2_2684(WX7785,WX7703,WX7728);
  and AND2_2685(WX7787,WX7702,WX7728);
  and AND2_2686(WX7789,WX7701,WX7728);
  and AND2_2687(WX7791,WX7700,WX7728);
  and AND2_2688(WX7793,WX7804,WX8761);
  and AND2_2689(WX7794,WX7800,WX7795);
  and AND2_2690(WX7797,CRC_OUT_3_31,WX8762);
  and AND2_2691(WX7798,WX10063,WX7799);
  and AND2_2692(WX7801,WX8243,WX8762);
  and AND2_2693(WX7802,WX8770,WX7803);
  and AND2_2694(WX7807,WX7818,WX8761);
  and AND2_2695(WX7808,WX7814,WX7809);
  and AND2_2696(WX7811,CRC_OUT_3_30,WX8762);
  and AND2_2697(WX7812,WX10070,WX7813);
  and AND2_2698(WX7815,WX8245,WX8762);
  and AND2_2699(WX7816,WX8777,WX7817);
  and AND2_2700(WX7821,WX7832,WX8761);
  and AND2_2701(WX7822,WX7828,WX7823);
  and AND2_2702(WX7825,CRC_OUT_3_29,WX8762);
  and AND2_2703(WX7826,WX10077,WX7827);
  and AND2_2704(WX7829,WX8247,WX8762);
  and AND2_2705(WX7830,WX8784,WX7831);
  and AND2_2706(WX7835,WX7846,WX8761);
  and AND2_2707(WX7836,WX7842,WX7837);
  and AND2_2708(WX7839,CRC_OUT_3_28,WX8762);
  and AND2_2709(WX7840,WX10084,WX7841);
  and AND2_2710(WX7843,WX8249,WX8762);
  and AND2_2711(WX7844,WX8791,WX7845);
  and AND2_2712(WX7849,WX7860,WX8761);
  and AND2_2713(WX7850,WX7856,WX7851);
  and AND2_2714(WX7853,CRC_OUT_3_27,WX8762);
  and AND2_2715(WX7854,WX10091,WX7855);
  and AND2_2716(WX7857,WX8251,WX8762);
  and AND2_2717(WX7858,WX8798,WX7859);
  and AND2_2718(WX7863,WX7874,WX8761);
  and AND2_2719(WX7864,WX7870,WX7865);
  and AND2_2720(WX7867,CRC_OUT_3_26,WX8762);
  and AND2_2721(WX7868,WX10098,WX7869);
  and AND2_2722(WX7871,WX8253,WX8762);
  and AND2_2723(WX7872,WX8805,WX7873);
  and AND2_2724(WX7877,WX7888,WX8761);
  and AND2_2725(WX7878,WX7884,WX7879);
  and AND2_2726(WX7881,CRC_OUT_3_25,WX8762);
  and AND2_2727(WX7882,WX10105,WX7883);
  and AND2_2728(WX7885,WX8255,WX8762);
  and AND2_2729(WX7886,WX8812,WX7887);
  and AND2_2730(WX7891,WX7902,WX8761);
  and AND2_2731(WX7892,WX7898,WX7893);
  and AND2_2732(WX7895,CRC_OUT_3_24,WX8762);
  and AND2_2733(WX7896,WX10112,WX7897);
  and AND2_2734(WX7899,WX8257,WX8762);
  and AND2_2735(WX7900,WX8819,WX7901);
  and AND2_2736(WX7905,WX7916,WX8761);
  and AND2_2737(WX7906,WX7912,WX7907);
  and AND2_2738(WX7909,CRC_OUT_3_23,WX8762);
  and AND2_2739(WX7910,WX10119,WX7911);
  and AND2_2740(WX7913,WX8259,WX8762);
  and AND2_2741(WX7914,WX8826,WX7915);
  and AND2_2742(WX7919,WX7930,WX8761);
  and AND2_2743(WX7920,WX7926,WX7921);
  and AND2_2744(WX7923,CRC_OUT_3_22,WX8762);
  and AND2_2745(WX7924,WX10126,WX7925);
  and AND2_2746(WX7927,WX8261,WX8762);
  and AND2_2747(WX7928,WX8833,WX7929);
  and AND2_2748(WX7933,WX7944,WX8761);
  and AND2_2749(WX7934,WX7940,WX7935);
  and AND2_2750(WX7937,CRC_OUT_3_21,WX8762);
  and AND2_2751(WX7938,WX10133,WX7939);
  and AND2_2752(WX7941,WX8263,WX8762);
  and AND2_2753(WX7942,WX8840,WX7943);
  and AND2_2754(WX7947,WX7958,WX8761);
  and AND2_2755(WX7948,WX7954,WX7949);
  and AND2_2756(WX7951,CRC_OUT_3_20,WX8762);
  and AND2_2757(WX7952,WX10140,WX7953);
  and AND2_2758(WX7955,WX8265,WX8762);
  and AND2_2759(WX7956,WX8847,WX7957);
  and AND2_2760(WX7961,WX7972,WX8761);
  and AND2_2761(WX7962,WX7968,WX7963);
  and AND2_2762(WX7965,CRC_OUT_3_19,WX8762);
  and AND2_2763(WX7966,WX10147,WX7967);
  and AND2_2764(WX7969,WX8267,WX8762);
  and AND2_2765(WX7970,WX8854,WX7971);
  and AND2_2766(WX7975,WX7986,WX8761);
  and AND2_2767(WX7976,WX7982,WX7977);
  and AND2_2768(WX7979,CRC_OUT_3_18,WX8762);
  and AND2_2769(WX7980,WX10154,WX7981);
  and AND2_2770(WX7983,WX8269,WX8762);
  and AND2_2771(WX7984,WX8861,WX7985);
  and AND2_2772(WX7989,WX8000,WX8761);
  and AND2_2773(WX7990,WX7996,WX7991);
  and AND2_2774(WX7993,CRC_OUT_3_17,WX8762);
  and AND2_2775(WX7994,WX10161,WX7995);
  and AND2_2776(WX7997,WX8271,WX8762);
  and AND2_2777(WX7998,WX8868,WX7999);
  and AND2_2778(WX8003,WX8014,WX8761);
  and AND2_2779(WX8004,WX8010,WX8005);
  and AND2_2780(WX8007,CRC_OUT_3_16,WX8762);
  and AND2_2781(WX8008,WX10168,WX8009);
  and AND2_2782(WX8011,WX8273,WX8762);
  and AND2_2783(WX8012,WX8875,WX8013);
  and AND2_2784(WX8017,WX8028,WX8761);
  and AND2_2785(WX8018,WX8024,WX8019);
  and AND2_2786(WX8021,CRC_OUT_3_15,WX8762);
  and AND2_2787(WX8022,WX10175,WX8023);
  and AND2_2788(WX8025,WX8275,WX8762);
  and AND2_2789(WX8026,WX8882,WX8027);
  and AND2_2790(WX8031,WX8042,WX8761);
  and AND2_2791(WX8032,WX8038,WX8033);
  and AND2_2792(WX8035,CRC_OUT_3_14,WX8762);
  and AND2_2793(WX8036,WX10182,WX8037);
  and AND2_2794(WX8039,WX8277,WX8762);
  and AND2_2795(WX8040,WX8889,WX8041);
  and AND2_2796(WX8045,WX8056,WX8761);
  and AND2_2797(WX8046,WX8052,WX8047);
  and AND2_2798(WX8049,CRC_OUT_3_13,WX8762);
  and AND2_2799(WX8050,WX10189,WX8051);
  and AND2_2800(WX8053,WX8279,WX8762);
  and AND2_2801(WX8054,WX8896,WX8055);
  and AND2_2802(WX8059,WX8070,WX8761);
  and AND2_2803(WX8060,WX8066,WX8061);
  and AND2_2804(WX8063,CRC_OUT_3_12,WX8762);
  and AND2_2805(WX8064,WX10196,WX8065);
  and AND2_2806(WX8067,WX8281,WX8762);
  and AND2_2807(WX8068,WX8903,WX8069);
  and AND2_2808(WX8073,WX8084,WX8761);
  and AND2_2809(WX8074,WX8080,WX8075);
  and AND2_2810(WX8077,CRC_OUT_3_11,WX8762);
  and AND2_2811(WX8078,WX10203,WX8079);
  and AND2_2812(WX8081,WX8283,WX8762);
  and AND2_2813(WX8082,WX8910,WX8083);
  and AND2_2814(WX8087,WX8098,WX8761);
  and AND2_2815(WX8088,WX8094,WX8089);
  and AND2_2816(WX8091,CRC_OUT_3_10,WX8762);
  and AND2_2817(WX8092,WX10210,WX8093);
  and AND2_2818(WX8095,WX8285,WX8762);
  and AND2_2819(WX8096,WX8917,WX8097);
  and AND2_2820(WX8101,WX8112,WX8761);
  and AND2_2821(WX8102,WX8108,WX8103);
  and AND2_2822(WX8105,CRC_OUT_3_9,WX8762);
  and AND2_2823(WX8106,WX10217,WX8107);
  and AND2_2824(WX8109,WX8287,WX8762);
  and AND2_2825(WX8110,WX8924,WX8111);
  and AND2_2826(WX8115,WX8126,WX8761);
  and AND2_2827(WX8116,WX8122,WX8117);
  and AND2_2828(WX8119,CRC_OUT_3_8,WX8762);
  and AND2_2829(WX8120,WX10224,WX8121);
  and AND2_2830(WX8123,WX8289,WX8762);
  and AND2_2831(WX8124,WX8931,WX8125);
  and AND2_2832(WX8129,WX8140,WX8761);
  and AND2_2833(WX8130,WX8136,WX8131);
  and AND2_2834(WX8133,CRC_OUT_3_7,WX8762);
  and AND2_2835(WX8134,WX10231,WX8135);
  and AND2_2836(WX8137,WX8291,WX8762);
  and AND2_2837(WX8138,WX8938,WX8139);
  and AND2_2838(WX8143,WX8154,WX8761);
  and AND2_2839(WX8144,WX8150,WX8145);
  and AND2_2840(WX8147,CRC_OUT_3_6,WX8762);
  and AND2_2841(WX8148,WX10238,WX8149);
  and AND2_2842(WX8151,WX8293,WX8762);
  and AND2_2843(WX8152,WX8945,WX8153);
  and AND2_2844(WX8157,WX8168,WX8761);
  and AND2_2845(WX8158,WX8164,WX8159);
  and AND2_2846(WX8161,CRC_OUT_3_5,WX8762);
  and AND2_2847(WX8162,WX10245,WX8163);
  and AND2_2848(WX8165,WX8295,WX8762);
  and AND2_2849(WX8166,WX8952,WX8167);
  and AND2_2850(WX8171,WX8182,WX8761);
  and AND2_2851(WX8172,WX8178,WX8173);
  and AND2_2852(WX8175,CRC_OUT_3_4,WX8762);
  and AND2_2853(WX8176,WX10252,WX8177);
  and AND2_2854(WX8179,WX8297,WX8762);
  and AND2_2855(WX8180,WX8959,WX8181);
  and AND2_2856(WX8185,WX8196,WX8761);
  and AND2_2857(WX8186,WX8192,WX8187);
  and AND2_2858(WX8189,CRC_OUT_3_3,WX8762);
  and AND2_2859(WX8190,WX10259,WX8191);
  and AND2_2860(WX8193,WX8299,WX8762);
  and AND2_2861(WX8194,WX8966,WX8195);
  and AND2_2862(WX8199,WX8210,WX8761);
  and AND2_2863(WX8200,WX8206,WX8201);
  and AND2_2864(WX8203,CRC_OUT_3_2,WX8762);
  and AND2_2865(WX8204,WX10266,WX8205);
  and AND2_2866(WX8207,WX8301,WX8762);
  and AND2_2867(WX8208,WX8973,WX8209);
  and AND2_2868(WX8213,WX8224,WX8761);
  and AND2_2869(WX8214,WX8220,WX8215);
  and AND2_2870(WX8217,CRC_OUT_3_1,WX8762);
  and AND2_2871(WX8218,WX10273,WX8219);
  and AND2_2872(WX8221,WX8303,WX8762);
  and AND2_2873(WX8222,WX8980,WX8223);
  and AND2_2874(WX8227,WX8238,WX8761);
  and AND2_2875(WX8228,WX8234,WX8229);
  and AND2_2876(WX8231,CRC_OUT_3_0,WX8762);
  and AND2_2877(WX8232,WX10280,WX8233);
  and AND2_2878(WX8235,WX8305,WX8762);
  and AND2_2879(WX8236,WX8987,WX8237);
  and AND2_2880(WX8242,WX8245,RESET);
  and AND2_2881(WX8244,WX8247,RESET);
  and AND2_2882(WX8246,WX8249,RESET);
  and AND2_2883(WX8248,WX8251,RESET);
  and AND2_2884(WX8250,WX8253,RESET);
  and AND2_2885(WX8252,WX8255,RESET);
  and AND2_2886(WX8254,WX8257,RESET);
  and AND2_2887(WX8256,WX8259,RESET);
  and AND2_2888(WX8258,WX8261,RESET);
  and AND2_2889(WX8260,WX8263,RESET);
  and AND2_2890(WX8262,WX8265,RESET);
  and AND2_2891(WX8264,WX8267,RESET);
  and AND2_2892(WX8266,WX8269,RESET);
  and AND2_2893(WX8268,WX8271,RESET);
  and AND2_2894(WX8270,WX8273,RESET);
  and AND2_2895(WX8272,WX8275,RESET);
  and AND2_2896(WX8274,WX8277,RESET);
  and AND2_2897(WX8276,WX8279,RESET);
  and AND2_2898(WX8278,WX8281,RESET);
  and AND2_2899(WX8280,WX8283,RESET);
  and AND2_2900(WX8282,WX8285,RESET);
  and AND2_2901(WX8284,WX8287,RESET);
  and AND2_2902(WX8286,WX8289,RESET);
  and AND2_2903(WX8288,WX8291,RESET);
  and AND2_2904(WX8290,WX8293,RESET);
  and AND2_2905(WX8292,WX8295,RESET);
  and AND2_2906(WX8294,WX8297,RESET);
  and AND2_2907(WX8296,WX8299,RESET);
  and AND2_2908(WX8298,WX8301,RESET);
  and AND2_2909(WX8300,WX8303,RESET);
  and AND2_2910(WX8302,WX8305,RESET);
  and AND2_2911(WX8304,WX8241,RESET);
  and AND2_2912(WX8402,WX7806,RESET);
  and AND2_2913(WX8404,WX7820,RESET);
  and AND2_2914(WX8406,WX7834,RESET);
  and AND2_2915(WX8408,WX7848,RESET);
  and AND2_2916(WX8410,WX7862,RESET);
  and AND2_2917(WX8412,WX7876,RESET);
  and AND2_2918(WX8414,WX7890,RESET);
  and AND2_2919(WX8416,WX7904,RESET);
  and AND2_2920(WX8418,WX7918,RESET);
  and AND2_2921(WX8420,WX7932,RESET);
  and AND2_2922(WX8422,WX7946,RESET);
  and AND2_2923(WX8424,WX7960,RESET);
  and AND2_2924(WX8426,WX7974,RESET);
  and AND2_2925(WX8428,WX7988,RESET);
  and AND2_2926(WX8430,WX8002,RESET);
  and AND2_2927(WX8432,WX8016,RESET);
  and AND2_2928(WX8434,WX8030,RESET);
  and AND2_2929(WX8436,WX8044,RESET);
  and AND2_2930(WX8438,WX8058,RESET);
  and AND2_2931(WX8440,WX8072,RESET);
  and AND2_2932(WX8442,WX8086,RESET);
  and AND2_2933(WX8444,WX8100,RESET);
  and AND2_2934(WX8446,WX8114,RESET);
  and AND2_2935(WX8448,WX8128,RESET);
  and AND2_2936(WX8450,WX8142,RESET);
  and AND2_2937(WX8452,WX8156,RESET);
  and AND2_2938(WX8454,WX8170,RESET);
  and AND2_2939(WX8456,WX8184,RESET);
  and AND2_2940(WX8458,WX8198,RESET);
  and AND2_2941(WX8460,WX8212,RESET);
  and AND2_2942(WX8462,WX8226,RESET);
  and AND2_2943(WX8464,WX8240,RESET);
  and AND2_2944(WX8466,WX8403,RESET);
  and AND2_2945(WX8468,WX8405,RESET);
  and AND2_2946(WX8470,WX8407,RESET);
  and AND2_2947(WX8472,WX8409,RESET);
  and AND2_2948(WX8474,WX8411,RESET);
  and AND2_2949(WX8476,WX8413,RESET);
  and AND2_2950(WX8478,WX8415,RESET);
  and AND2_2951(WX8480,WX8417,RESET);
  and AND2_2952(WX8482,WX8419,RESET);
  and AND2_2953(WX8484,WX8421,RESET);
  and AND2_2954(WX8486,WX8423,RESET);
  and AND2_2955(WX8488,WX8425,RESET);
  and AND2_2956(WX8490,WX8427,RESET);
  and AND2_2957(WX8492,WX8429,RESET);
  and AND2_2958(WX8494,WX8431,RESET);
  and AND2_2959(WX8496,WX8433,RESET);
  and AND2_2960(WX8498,WX8435,RESET);
  and AND2_2961(WX8500,WX8437,RESET);
  and AND2_2962(WX8502,WX8439,RESET);
  and AND2_2963(WX8504,WX8441,RESET);
  and AND2_2964(WX8506,WX8443,RESET);
  and AND2_2965(WX8508,WX8445,RESET);
  and AND2_2966(WX8510,WX8447,RESET);
  and AND2_2967(WX8512,WX8449,RESET);
  and AND2_2968(WX8514,WX8451,RESET);
  and AND2_2969(WX8516,WX8453,RESET);
  and AND2_2970(WX8518,WX8455,RESET);
  and AND2_2971(WX8520,WX8457,RESET);
  and AND2_2972(WX8522,WX8459,RESET);
  and AND2_2973(WX8524,WX8461,RESET);
  and AND2_2974(WX8526,WX8463,RESET);
  and AND2_2975(WX8528,WX8465,RESET);
  and AND2_2976(WX8530,WX8467,RESET);
  and AND2_2977(WX8532,WX8469,RESET);
  and AND2_2978(WX8534,WX8471,RESET);
  and AND2_2979(WX8536,WX8473,RESET);
  and AND2_2980(WX8538,WX8475,RESET);
  and AND2_2981(WX8540,WX8477,RESET);
  and AND2_2982(WX8542,WX8479,RESET);
  and AND2_2983(WX8544,WX8481,RESET);
  and AND2_2984(WX8546,WX8483,RESET);
  and AND2_2985(WX8548,WX8485,RESET);
  and AND2_2986(WX8550,WX8487,RESET);
  and AND2_2987(WX8552,WX8489,RESET);
  and AND2_2988(WX8554,WX8491,RESET);
  and AND2_2989(WX8556,WX8493,RESET);
  and AND2_2990(WX8558,WX8495,RESET);
  and AND2_2991(WX8560,WX8497,RESET);
  and AND2_2992(WX8562,WX8499,RESET);
  and AND2_2993(WX8564,WX8501,RESET);
  and AND2_2994(WX8566,WX8503,RESET);
  and AND2_2995(WX8568,WX8505,RESET);
  and AND2_2996(WX8570,WX8507,RESET);
  and AND2_2997(WX8572,WX8509,RESET);
  and AND2_2998(WX8574,WX8511,RESET);
  and AND2_2999(WX8576,WX8513,RESET);
  and AND2_3000(WX8578,WX8515,RESET);
  and AND2_3001(WX8580,WX8517,RESET);
  and AND2_3002(WX8582,WX8519,RESET);
  and AND2_3003(WX8584,WX8521,RESET);
  and AND2_3004(WX8586,WX8523,RESET);
  and AND2_3005(WX8588,WX8525,RESET);
  and AND2_3006(WX8590,WX8527,RESET);
  and AND2_3007(WX8592,WX8529,RESET);
  and AND2_3008(WX8594,WX8531,RESET);
  and AND2_3009(WX8596,WX8533,RESET);
  and AND2_3010(WX8598,WX8535,RESET);
  and AND2_3011(WX8600,WX8537,RESET);
  and AND2_3012(WX8602,WX8539,RESET);
  and AND2_3013(WX8604,WX8541,RESET);
  and AND2_3014(WX8606,WX8543,RESET);
  and AND2_3015(WX8608,WX8545,RESET);
  and AND2_3016(WX8610,WX8547,RESET);
  and AND2_3017(WX8612,WX8549,RESET);
  and AND2_3018(WX8614,WX8551,RESET);
  and AND2_3019(WX8616,WX8553,RESET);
  and AND2_3020(WX8618,WX8555,RESET);
  and AND2_3021(WX8620,WX8557,RESET);
  and AND2_3022(WX8622,WX8559,RESET);
  and AND2_3023(WX8624,WX8561,RESET);
  and AND2_3024(WX8626,WX8563,RESET);
  and AND2_3025(WX8628,WX8565,RESET);
  and AND2_3026(WX8630,WX8567,RESET);
  and AND2_3027(WX8632,WX8569,RESET);
  and AND2_3028(WX8634,WX8571,RESET);
  and AND2_3029(WX8636,WX8573,RESET);
  and AND2_3030(WX8638,WX8575,RESET);
  and AND2_3031(WX8640,WX8577,RESET);
  and AND2_3032(WX8642,WX8579,RESET);
  and AND2_3033(WX8644,WX8581,RESET);
  and AND2_3034(WX8646,WX8583,RESET);
  and AND2_3035(WX8648,WX8585,RESET);
  and AND2_3036(WX8650,WX8587,RESET);
  and AND2_3037(WX8652,WX8589,RESET);
  and AND2_3038(WX8654,WX8591,RESET);
  and AND2_3039(WX8656,WX8593,RESET);
  and AND2_3040(WX8765,WX8764,WX8763);
  and AND2_3041(WX8766,WX8338,WX8767);
  and AND2_3042(WX8772,WX8771,WX8763);
  and AND2_3043(WX8773,WX8339,WX8774);
  and AND2_3044(WX8779,WX8778,WX8763);
  and AND2_3045(WX8780,WX8340,WX8781);
  and AND2_3046(WX8786,WX8785,WX8763);
  and AND2_3047(WX8787,WX8341,WX8788);
  and AND2_3048(WX8793,WX8792,WX8763);
  and AND2_3049(WX8794,WX8342,WX8795);
  and AND2_3050(WX8800,WX8799,WX8763);
  and AND2_3051(WX8801,WX8343,WX8802);
  and AND2_3052(WX8807,WX8806,WX8763);
  and AND2_3053(WX8808,WX8344,WX8809);
  and AND2_3054(WX8814,WX8813,WX8763);
  and AND2_3055(WX8815,WX8345,WX8816);
  and AND2_3056(WX8821,WX8820,WX8763);
  and AND2_3057(WX8822,WX8346,WX8823);
  and AND2_3058(WX8828,WX8827,WX8763);
  and AND2_3059(WX8829,WX8347,WX8830);
  and AND2_3060(WX8835,WX8834,WX8763);
  and AND2_3061(WX8836,WX8348,WX8837);
  and AND2_3062(WX8842,WX8841,WX8763);
  and AND2_3063(WX8843,WX8349,WX8844);
  and AND2_3064(WX8849,WX8848,WX8763);
  and AND2_3065(WX8850,WX8350,WX8851);
  and AND2_3066(WX8856,WX8855,WX8763);
  and AND2_3067(WX8857,WX8351,WX8858);
  and AND2_3068(WX8863,WX8862,WX8763);
  and AND2_3069(WX8864,WX8352,WX8865);
  and AND2_3070(WX8870,WX8869,WX8763);
  and AND2_3071(WX8871,WX8353,WX8872);
  and AND2_3072(WX8877,WX8876,WX8763);
  and AND2_3073(WX8878,WX8354,WX8879);
  and AND2_3074(WX8884,WX8883,WX8763);
  and AND2_3075(WX8885,WX8355,WX8886);
  and AND2_3076(WX8891,WX8890,WX8763);
  and AND2_3077(WX8892,WX8356,WX8893);
  and AND2_3078(WX8898,WX8897,WX8763);
  and AND2_3079(WX8899,WX8357,WX8900);
  and AND2_3080(WX8905,WX8904,WX8763);
  and AND2_3081(WX8906,WX8358,WX8907);
  and AND2_3082(WX8912,WX8911,WX8763);
  and AND2_3083(WX8913,WX8359,WX8914);
  and AND2_3084(WX8919,WX8918,WX8763);
  and AND2_3085(WX8920,WX8360,WX8921);
  and AND2_3086(WX8926,WX8925,WX8763);
  and AND2_3087(WX8927,WX8361,WX8928);
  and AND2_3088(WX8933,WX8932,WX8763);
  and AND2_3089(WX8934,WX8362,WX8935);
  and AND2_3090(WX8940,WX8939,WX8763);
  and AND2_3091(WX8941,WX8363,WX8942);
  and AND2_3092(WX8947,WX8946,WX8763);
  and AND2_3093(WX8948,WX8364,WX8949);
  and AND2_3094(WX8954,WX8953,WX8763);
  and AND2_3095(WX8955,WX8365,WX8956);
  and AND2_3096(WX8961,WX8960,WX8763);
  and AND2_3097(WX8962,WX8366,WX8963);
  and AND2_3098(WX8968,WX8967,WX8763);
  and AND2_3099(WX8969,WX8367,WX8970);
  and AND2_3100(WX8975,WX8974,WX8763);
  and AND2_3101(WX8976,WX8368,WX8977);
  and AND2_3102(WX8982,WX8981,WX8763);
  and AND2_3103(WX8983,WX8369,WX8984);
  and AND2_3104(WX9022,WX8992,WX9021);
  and AND2_3105(WX9024,WX9020,WX9021);
  and AND2_3106(WX9026,WX9019,WX9021);
  and AND2_3107(WX9028,WX9018,WX9021);
  and AND2_3108(WX9030,WX8991,WX9021);
  and AND2_3109(WX9032,WX9017,WX9021);
  and AND2_3110(WX9034,WX9016,WX9021);
  and AND2_3111(WX9036,WX9015,WX9021);
  and AND2_3112(WX9038,WX9014,WX9021);
  and AND2_3113(WX9040,WX9013,WX9021);
  and AND2_3114(WX9042,WX9012,WX9021);
  and AND2_3115(WX9044,WX8990,WX9021);
  and AND2_3116(WX9046,WX9011,WX9021);
  and AND2_3117(WX9048,WX9010,WX9021);
  and AND2_3118(WX9050,WX9009,WX9021);
  and AND2_3119(WX9052,WX9008,WX9021);
  and AND2_3120(WX9054,WX8989,WX9021);
  and AND2_3121(WX9056,WX9007,WX9021);
  and AND2_3122(WX9058,WX9006,WX9021);
  and AND2_3123(WX9060,WX9005,WX9021);
  and AND2_3124(WX9062,WX9004,WX9021);
  and AND2_3125(WX9064,WX9003,WX9021);
  and AND2_3126(WX9066,WX9002,WX9021);
  and AND2_3127(WX9068,WX9001,WX9021);
  and AND2_3128(WX9070,WX9000,WX9021);
  and AND2_3129(WX9072,WX8999,WX9021);
  and AND2_3130(WX9074,WX8998,WX9021);
  and AND2_3131(WX9076,WX8997,WX9021);
  and AND2_3132(WX9078,WX8996,WX9021);
  and AND2_3133(WX9080,WX8995,WX9021);
  and AND2_3134(WX9082,WX8994,WX9021);
  and AND2_3135(WX9084,WX8993,WX9021);
  and AND2_3136(WX9086,WX9097,WX10054);
  and AND2_3137(WX9087,WX9093,WX9088);
  and AND2_3138(WX9090,CRC_OUT_2_31,WX10055);
  and AND2_3139(WX9091,WX11356,WX9092);
  and AND2_3140(WX9094,WX9536,WX10055);
  and AND2_3141(WX9095,WX10063,WX9096);
  and AND2_3142(WX9100,WX9111,WX10054);
  and AND2_3143(WX9101,WX9107,WX9102);
  and AND2_3144(WX9104,CRC_OUT_2_30,WX10055);
  and AND2_3145(WX9105,WX11363,WX9106);
  and AND2_3146(WX9108,WX9538,WX10055);
  and AND2_3147(WX9109,WX10070,WX9110);
  and AND2_3148(WX9114,WX9125,WX10054);
  and AND2_3149(WX9115,WX9121,WX9116);
  and AND2_3150(WX9118,CRC_OUT_2_29,WX10055);
  and AND2_3151(WX9119,WX11370,WX9120);
  and AND2_3152(WX9122,WX9540,WX10055);
  and AND2_3153(WX9123,WX10077,WX9124);
  and AND2_3154(WX9128,WX9139,WX10054);
  and AND2_3155(WX9129,WX9135,WX9130);
  and AND2_3156(WX9132,CRC_OUT_2_28,WX10055);
  and AND2_3157(WX9133,WX11377,WX9134);
  and AND2_3158(WX9136,WX9542,WX10055);
  and AND2_3159(WX9137,WX10084,WX9138);
  and AND2_3160(WX9142,WX9153,WX10054);
  and AND2_3161(WX9143,WX9149,WX9144);
  and AND2_3162(WX9146,CRC_OUT_2_27,WX10055);
  and AND2_3163(WX9147,WX11384,WX9148);
  and AND2_3164(WX9150,WX9544,WX10055);
  and AND2_3165(WX9151,WX10091,WX9152);
  and AND2_3166(WX9156,WX9167,WX10054);
  and AND2_3167(WX9157,WX9163,WX9158);
  and AND2_3168(WX9160,CRC_OUT_2_26,WX10055);
  and AND2_3169(WX9161,WX11391,WX9162);
  and AND2_3170(WX9164,WX9546,WX10055);
  and AND2_3171(WX9165,WX10098,WX9166);
  and AND2_3172(WX9170,WX9181,WX10054);
  and AND2_3173(WX9171,WX9177,WX9172);
  and AND2_3174(WX9174,CRC_OUT_2_25,WX10055);
  and AND2_3175(WX9175,WX11398,WX9176);
  and AND2_3176(WX9178,WX9548,WX10055);
  and AND2_3177(WX9179,WX10105,WX9180);
  and AND2_3178(WX9184,WX9195,WX10054);
  and AND2_3179(WX9185,WX9191,WX9186);
  and AND2_3180(WX9188,CRC_OUT_2_24,WX10055);
  and AND2_3181(WX9189,WX11405,WX9190);
  and AND2_3182(WX9192,WX9550,WX10055);
  and AND2_3183(WX9193,WX10112,WX9194);
  and AND2_3184(WX9198,WX9209,WX10054);
  and AND2_3185(WX9199,WX9205,WX9200);
  and AND2_3186(WX9202,CRC_OUT_2_23,WX10055);
  and AND2_3187(WX9203,WX11412,WX9204);
  and AND2_3188(WX9206,WX9552,WX10055);
  and AND2_3189(WX9207,WX10119,WX9208);
  and AND2_3190(WX9212,WX9223,WX10054);
  and AND2_3191(WX9213,WX9219,WX9214);
  and AND2_3192(WX9216,CRC_OUT_2_22,WX10055);
  and AND2_3193(WX9217,WX11419,WX9218);
  and AND2_3194(WX9220,WX9554,WX10055);
  and AND2_3195(WX9221,WX10126,WX9222);
  and AND2_3196(WX9226,WX9237,WX10054);
  and AND2_3197(WX9227,WX9233,WX9228);
  and AND2_3198(WX9230,CRC_OUT_2_21,WX10055);
  and AND2_3199(WX9231,WX11426,WX9232);
  and AND2_3200(WX9234,WX9556,WX10055);
  and AND2_3201(WX9235,WX10133,WX9236);
  and AND2_3202(WX9240,WX9251,WX10054);
  and AND2_3203(WX9241,WX9247,WX9242);
  and AND2_3204(WX9244,CRC_OUT_2_20,WX10055);
  and AND2_3205(WX9245,WX11433,WX9246);
  and AND2_3206(WX9248,WX9558,WX10055);
  and AND2_3207(WX9249,WX10140,WX9250);
  and AND2_3208(WX9254,WX9265,WX10054);
  and AND2_3209(WX9255,WX9261,WX9256);
  and AND2_3210(WX9258,CRC_OUT_2_19,WX10055);
  and AND2_3211(WX9259,WX11440,WX9260);
  and AND2_3212(WX9262,WX9560,WX10055);
  and AND2_3213(WX9263,WX10147,WX9264);
  and AND2_3214(WX9268,WX9279,WX10054);
  and AND2_3215(WX9269,WX9275,WX9270);
  and AND2_3216(WX9272,CRC_OUT_2_18,WX10055);
  and AND2_3217(WX9273,WX11447,WX9274);
  and AND2_3218(WX9276,WX9562,WX10055);
  and AND2_3219(WX9277,WX10154,WX9278);
  and AND2_3220(WX9282,WX9293,WX10054);
  and AND2_3221(WX9283,WX9289,WX9284);
  and AND2_3222(WX9286,CRC_OUT_2_17,WX10055);
  and AND2_3223(WX9287,WX11454,WX9288);
  and AND2_3224(WX9290,WX9564,WX10055);
  and AND2_3225(WX9291,WX10161,WX9292);
  and AND2_3226(WX9296,WX9307,WX10054);
  and AND2_3227(WX9297,WX9303,WX9298);
  and AND2_3228(WX9300,CRC_OUT_2_16,WX10055);
  and AND2_3229(WX9301,WX11461,WX9302);
  and AND2_3230(WX9304,WX9566,WX10055);
  and AND2_3231(WX9305,WX10168,WX9306);
  and AND2_3232(WX9310,WX9321,WX10054);
  and AND2_3233(WX9311,WX9317,WX9312);
  and AND2_3234(WX9314,CRC_OUT_2_15,WX10055);
  and AND2_3235(WX9315,WX11468,WX9316);
  and AND2_3236(WX9318,WX9568,WX10055);
  and AND2_3237(WX9319,WX10175,WX9320);
  and AND2_3238(WX9324,WX9335,WX10054);
  and AND2_3239(WX9325,WX9331,WX9326);
  and AND2_3240(WX9328,CRC_OUT_2_14,WX10055);
  and AND2_3241(WX9329,WX11475,WX9330);
  and AND2_3242(WX9332,WX9570,WX10055);
  and AND2_3243(WX9333,WX10182,WX9334);
  and AND2_3244(WX9338,WX9349,WX10054);
  and AND2_3245(WX9339,WX9345,WX9340);
  and AND2_3246(WX9342,CRC_OUT_2_13,WX10055);
  and AND2_3247(WX9343,WX11482,WX9344);
  and AND2_3248(WX9346,WX9572,WX10055);
  and AND2_3249(WX9347,WX10189,WX9348);
  and AND2_3250(WX9352,WX9363,WX10054);
  and AND2_3251(WX9353,WX9359,WX9354);
  and AND2_3252(WX9356,CRC_OUT_2_12,WX10055);
  and AND2_3253(WX9357,WX11489,WX9358);
  and AND2_3254(WX9360,WX9574,WX10055);
  and AND2_3255(WX9361,WX10196,WX9362);
  and AND2_3256(WX9366,WX9377,WX10054);
  and AND2_3257(WX9367,WX9373,WX9368);
  and AND2_3258(WX9370,CRC_OUT_2_11,WX10055);
  and AND2_3259(WX9371,WX11496,WX9372);
  and AND2_3260(WX9374,WX9576,WX10055);
  and AND2_3261(WX9375,WX10203,WX9376);
  and AND2_3262(WX9380,WX9391,WX10054);
  and AND2_3263(WX9381,WX9387,WX9382);
  and AND2_3264(WX9384,CRC_OUT_2_10,WX10055);
  and AND2_3265(WX9385,WX11503,WX9386);
  and AND2_3266(WX9388,WX9578,WX10055);
  and AND2_3267(WX9389,WX10210,WX9390);
  and AND2_3268(WX9394,WX9405,WX10054);
  and AND2_3269(WX9395,WX9401,WX9396);
  and AND2_3270(WX9398,CRC_OUT_2_9,WX10055);
  and AND2_3271(WX9399,WX11510,WX9400);
  and AND2_3272(WX9402,WX9580,WX10055);
  and AND2_3273(WX9403,WX10217,WX9404);
  and AND2_3274(WX9408,WX9419,WX10054);
  and AND2_3275(WX9409,WX9415,WX9410);
  and AND2_3276(WX9412,CRC_OUT_2_8,WX10055);
  and AND2_3277(WX9413,WX11517,WX9414);
  and AND2_3278(WX9416,WX9582,WX10055);
  and AND2_3279(WX9417,WX10224,WX9418);
  and AND2_3280(WX9422,WX9433,WX10054);
  and AND2_3281(WX9423,WX9429,WX9424);
  and AND2_3282(WX9426,CRC_OUT_2_7,WX10055);
  and AND2_3283(WX9427,WX11524,WX9428);
  and AND2_3284(WX9430,WX9584,WX10055);
  and AND2_3285(WX9431,WX10231,WX9432);
  and AND2_3286(WX9436,WX9447,WX10054);
  and AND2_3287(WX9437,WX9443,WX9438);
  and AND2_3288(WX9440,CRC_OUT_2_6,WX10055);
  and AND2_3289(WX9441,WX11531,WX9442);
  and AND2_3290(WX9444,WX9586,WX10055);
  and AND2_3291(WX9445,WX10238,WX9446);
  and AND2_3292(WX9450,WX9461,WX10054);
  and AND2_3293(WX9451,WX9457,WX9452);
  and AND2_3294(WX9454,CRC_OUT_2_5,WX10055);
  and AND2_3295(WX9455,WX11538,WX9456);
  and AND2_3296(WX9458,WX9588,WX10055);
  and AND2_3297(WX9459,WX10245,WX9460);
  and AND2_3298(WX9464,WX9475,WX10054);
  and AND2_3299(WX9465,WX9471,WX9466);
  and AND2_3300(WX9468,CRC_OUT_2_4,WX10055);
  and AND2_3301(WX9469,WX11545,WX9470);
  and AND2_3302(WX9472,WX9590,WX10055);
  and AND2_3303(WX9473,WX10252,WX9474);
  and AND2_3304(WX9478,WX9489,WX10054);
  and AND2_3305(WX9479,WX9485,WX9480);
  and AND2_3306(WX9482,CRC_OUT_2_3,WX10055);
  and AND2_3307(WX9483,WX11552,WX9484);
  and AND2_3308(WX9486,WX9592,WX10055);
  and AND2_3309(WX9487,WX10259,WX9488);
  and AND2_3310(WX9492,WX9503,WX10054);
  and AND2_3311(WX9493,WX9499,WX9494);
  and AND2_3312(WX9496,CRC_OUT_2_2,WX10055);
  and AND2_3313(WX9497,WX11559,WX9498);
  and AND2_3314(WX9500,WX9594,WX10055);
  and AND2_3315(WX9501,WX10266,WX9502);
  and AND2_3316(WX9506,WX9517,WX10054);
  and AND2_3317(WX9507,WX9513,WX9508);
  and AND2_3318(WX9510,CRC_OUT_2_1,WX10055);
  and AND2_3319(WX9511,WX11566,WX9512);
  and AND2_3320(WX9514,WX9596,WX10055);
  and AND2_3321(WX9515,WX10273,WX9516);
  and AND2_3322(WX9520,WX9531,WX10054);
  and AND2_3323(WX9521,WX9527,WX9522);
  and AND2_3324(WX9524,CRC_OUT_2_0,WX10055);
  and AND2_3325(WX9525,WX11573,WX9526);
  and AND2_3326(WX9528,WX9598,WX10055);
  and AND2_3327(WX9529,WX10280,WX9530);
  and AND2_3328(WX9535,WX9538,RESET);
  and AND2_3329(WX9537,WX9540,RESET);
  and AND2_3330(WX9539,WX9542,RESET);
  and AND2_3331(WX9541,WX9544,RESET);
  and AND2_3332(WX9543,WX9546,RESET);
  and AND2_3333(WX9545,WX9548,RESET);
  and AND2_3334(WX9547,WX9550,RESET);
  and AND2_3335(WX9549,WX9552,RESET);
  and AND2_3336(WX9551,WX9554,RESET);
  and AND2_3337(WX9553,WX9556,RESET);
  and AND2_3338(WX9555,WX9558,RESET);
  and AND2_3339(WX9557,WX9560,RESET);
  and AND2_3340(WX9559,WX9562,RESET);
  and AND2_3341(WX9561,WX9564,RESET);
  and AND2_3342(WX9563,WX9566,RESET);
  and AND2_3343(WX9565,WX9568,RESET);
  and AND2_3344(WX9567,WX9570,RESET);
  and AND2_3345(WX9569,WX9572,RESET);
  and AND2_3346(WX9571,WX9574,RESET);
  and AND2_3347(WX9573,WX9576,RESET);
  and AND2_3348(WX9575,WX9578,RESET);
  and AND2_3349(WX9577,WX9580,RESET);
  and AND2_3350(WX9579,WX9582,RESET);
  and AND2_3351(WX9581,WX9584,RESET);
  and AND2_3352(WX9583,WX9586,RESET);
  and AND2_3353(WX9585,WX9588,RESET);
  and AND2_3354(WX9587,WX9590,RESET);
  and AND2_3355(WX9589,WX9592,RESET);
  and AND2_3356(WX9591,WX9594,RESET);
  and AND2_3357(WX9593,WX9596,RESET);
  and AND2_3358(WX9595,WX9598,RESET);
  and AND2_3359(WX9597,WX9534,RESET);
  and AND2_3360(WX9695,WX9099,RESET);
  and AND2_3361(WX9697,WX9113,RESET);
  and AND2_3362(WX9699,WX9127,RESET);
  and AND2_3363(WX9701,WX9141,RESET);
  and AND2_3364(WX9703,WX9155,RESET);
  and AND2_3365(WX9705,WX9169,RESET);
  and AND2_3366(WX9707,WX9183,RESET);
  and AND2_3367(WX9709,WX9197,RESET);
  and AND2_3368(WX9711,WX9211,RESET);
  and AND2_3369(WX9713,WX9225,RESET);
  and AND2_3370(WX9715,WX9239,RESET);
  and AND2_3371(WX9717,WX9253,RESET);
  and AND2_3372(WX9719,WX9267,RESET);
  and AND2_3373(WX9721,WX9281,RESET);
  and AND2_3374(WX9723,WX9295,RESET);
  and AND2_3375(WX9725,WX9309,RESET);
  and AND2_3376(WX9727,WX9323,RESET);
  and AND2_3377(WX9729,WX9337,RESET);
  and AND2_3378(WX9731,WX9351,RESET);
  and AND2_3379(WX9733,WX9365,RESET);
  and AND2_3380(WX9735,WX9379,RESET);
  and AND2_3381(WX9737,WX9393,RESET);
  and AND2_3382(WX9739,WX9407,RESET);
  and AND2_3383(WX9741,WX9421,RESET);
  and AND2_3384(WX9743,WX9435,RESET);
  and AND2_3385(WX9745,WX9449,RESET);
  and AND2_3386(WX9747,WX9463,RESET);
  and AND2_3387(WX9749,WX9477,RESET);
  and AND2_3388(WX9751,WX9491,RESET);
  and AND2_3389(WX9753,WX9505,RESET);
  and AND2_3390(WX9755,WX9519,RESET);
  and AND2_3391(WX9757,WX9533,RESET);
  and AND2_3392(WX9759,WX9696,RESET);
  and AND2_3393(WX9761,WX9698,RESET);
  and AND2_3394(WX9763,WX9700,RESET);
  and AND2_3395(WX9765,WX9702,RESET);
  and AND2_3396(WX9767,WX9704,RESET);
  and AND2_3397(WX9769,WX9706,RESET);
  and AND2_3398(WX9771,WX9708,RESET);
  and AND2_3399(WX9773,WX9710,RESET);
  and AND2_3400(WX9775,WX9712,RESET);
  and AND2_3401(WX9777,WX9714,RESET);
  and AND2_3402(WX9779,WX9716,RESET);
  and AND2_3403(WX9781,WX9718,RESET);
  and AND2_3404(WX9783,WX9720,RESET);
  and AND2_3405(WX9785,WX9722,RESET);
  and AND2_3406(WX9787,WX9724,RESET);
  and AND2_3407(WX9789,WX9726,RESET);
  and AND2_3408(WX9791,WX9728,RESET);
  and AND2_3409(WX9793,WX9730,RESET);
  and AND2_3410(WX9795,WX9732,RESET);
  and AND2_3411(WX9797,WX9734,RESET);
  and AND2_3412(WX9799,WX9736,RESET);
  and AND2_3413(WX9801,WX9738,RESET);
  and AND2_3414(WX9803,WX9740,RESET);
  and AND2_3415(WX9805,WX9742,RESET);
  and AND2_3416(WX9807,WX9744,RESET);
  and AND2_3417(WX9809,WX9746,RESET);
  and AND2_3418(WX9811,WX9748,RESET);
  and AND2_3419(WX9813,WX9750,RESET);
  and AND2_3420(WX9815,WX9752,RESET);
  and AND2_3421(WX9817,WX9754,RESET);
  and AND2_3422(WX9819,WX9756,RESET);
  and AND2_3423(WX9821,WX9758,RESET);
  and AND2_3424(WX9823,WX9760,RESET);
  and AND2_3425(WX9825,WX9762,RESET);
  and AND2_3426(WX9827,WX9764,RESET);
  and AND2_3427(WX9829,WX9766,RESET);
  and AND2_3428(WX9831,WX9768,RESET);
  and AND2_3429(WX9833,WX9770,RESET);
  and AND2_3430(WX9835,WX9772,RESET);
  and AND2_3431(WX9837,WX9774,RESET);
  and AND2_3432(WX9839,WX9776,RESET);
  and AND2_3433(WX9841,WX9778,RESET);
  and AND2_3434(WX9843,WX9780,RESET);
  and AND2_3435(WX9845,WX9782,RESET);
  and AND2_3436(WX9847,WX9784,RESET);
  and AND2_3437(WX9849,WX9786,RESET);
  and AND2_3438(WX9851,WX9788,RESET);
  and AND2_3439(WX9853,WX9790,RESET);
  and AND2_3440(WX9855,WX9792,RESET);
  and AND2_3441(WX9857,WX9794,RESET);
  and AND2_3442(WX9859,WX9796,RESET);
  and AND2_3443(WX9861,WX9798,RESET);
  and AND2_3444(WX9863,WX9800,RESET);
  and AND2_3445(WX9865,WX9802,RESET);
  and AND2_3446(WX9867,WX9804,RESET);
  and AND2_3447(WX9869,WX9806,RESET);
  and AND2_3448(WX9871,WX9808,RESET);
  and AND2_3449(WX9873,WX9810,RESET);
  and AND2_3450(WX9875,WX9812,RESET);
  and AND2_3451(WX9877,WX9814,RESET);
  and AND2_3452(WX9879,WX9816,RESET);
  and AND2_3453(WX9881,WX9818,RESET);
  and AND2_3454(WX9883,WX9820,RESET);
  and AND2_3455(WX9885,WX9822,RESET);
  and AND2_3456(WX9887,WX9824,RESET);
  and AND2_3457(WX9889,WX9826,RESET);
  and AND2_3458(WX9891,WX9828,RESET);
  and AND2_3459(WX9893,WX9830,RESET);
  and AND2_3460(WX9895,WX9832,RESET);
  and AND2_3461(WX9897,WX9834,RESET);
  and AND2_3462(WX9899,WX9836,RESET);
  and AND2_3463(WX9901,WX9838,RESET);
  and AND2_3464(WX9903,WX9840,RESET);
  and AND2_3465(WX9905,WX9842,RESET);
  and AND2_3466(WX9907,WX9844,RESET);
  and AND2_3467(WX9909,WX9846,RESET);
  and AND2_3468(WX9911,WX9848,RESET);
  and AND2_3469(WX9913,WX9850,RESET);
  and AND2_3470(WX9915,WX9852,RESET);
  and AND2_3471(WX9917,WX9854,RESET);
  and AND2_3472(WX9919,WX9856,RESET);
  and AND2_3473(WX9921,WX9858,RESET);
  and AND2_3474(WX9923,WX9860,RESET);
  and AND2_3475(WX9925,WX9862,RESET);
  and AND2_3476(WX9927,WX9864,RESET);
  and AND2_3477(WX9929,WX9866,RESET);
  and AND2_3478(WX9931,WX9868,RESET);
  and AND2_3479(WX9933,WX9870,RESET);
  and AND2_3480(WX9935,WX9872,RESET);
  and AND2_3481(WX9937,WX9874,RESET);
  and AND2_3482(WX9939,WX9876,RESET);
  and AND2_3483(WX9941,WX9878,RESET);
  and AND2_3484(WX9943,WX9880,RESET);
  and AND2_3485(WX9945,WX9882,RESET);
  and AND2_3486(WX9947,WX9884,RESET);
  and AND2_3487(WX9949,WX9886,RESET);
  and AND2_3488(WX10058,WX10057,WX10056);
  and AND2_3489(WX10059,WX9631,WX10060);
  and AND2_3490(WX10065,WX10064,WX10056);
  and AND2_3491(WX10066,WX9632,WX10067);
  and AND2_3492(WX10072,WX10071,WX10056);
  and AND2_3493(WX10073,WX9633,WX10074);
  and AND2_3494(WX10079,WX10078,WX10056);
  and AND2_3495(WX10080,WX9634,WX10081);
  and AND2_3496(WX10086,WX10085,WX10056);
  and AND2_3497(WX10087,WX9635,WX10088);
  and AND2_3498(WX10093,WX10092,WX10056);
  and AND2_3499(WX10094,WX9636,WX10095);
  and AND2_3500(WX10100,WX10099,WX10056);
  and AND2_3501(WX10101,WX9637,WX10102);
  and AND2_3502(WX10107,WX10106,WX10056);
  and AND2_3503(WX10108,WX9638,WX10109);
  and AND2_3504(WX10114,WX10113,WX10056);
  and AND2_3505(WX10115,WX9639,WX10116);
  and AND2_3506(WX10121,WX10120,WX10056);
  and AND2_3507(WX10122,WX9640,WX10123);
  and AND2_3508(WX10128,WX10127,WX10056);
  and AND2_3509(WX10129,WX9641,WX10130);
  and AND2_3510(WX10135,WX10134,WX10056);
  and AND2_3511(WX10136,WX9642,WX10137);
  and AND2_3512(WX10142,WX10141,WX10056);
  and AND2_3513(WX10143,WX9643,WX10144);
  and AND2_3514(WX10149,WX10148,WX10056);
  and AND2_3515(WX10150,WX9644,WX10151);
  and AND2_3516(WX10156,WX10155,WX10056);
  and AND2_3517(WX10157,WX9645,WX10158);
  and AND2_3518(WX10163,WX10162,WX10056);
  and AND2_3519(WX10164,WX9646,WX10165);
  and AND2_3520(WX10170,WX10169,WX10056);
  and AND2_3521(WX10171,WX9647,WX10172);
  and AND2_3522(WX10177,WX10176,WX10056);
  and AND2_3523(WX10178,WX9648,WX10179);
  and AND2_3524(WX10184,WX10183,WX10056);
  and AND2_3525(WX10185,WX9649,WX10186);
  and AND2_3526(WX10191,WX10190,WX10056);
  and AND2_3527(WX10192,WX9650,WX10193);
  and AND2_3528(WX10198,WX10197,WX10056);
  and AND2_3529(WX10199,WX9651,WX10200);
  and AND2_3530(WX10205,WX10204,WX10056);
  and AND2_3531(WX10206,WX9652,WX10207);
  and AND2_3532(WX10212,WX10211,WX10056);
  and AND2_3533(WX10213,WX9653,WX10214);
  and AND2_3534(WX10219,WX10218,WX10056);
  and AND2_3535(WX10220,WX9654,WX10221);
  and AND2_3536(WX10226,WX10225,WX10056);
  and AND2_3537(WX10227,WX9655,WX10228);
  and AND2_3538(WX10233,WX10232,WX10056);
  and AND2_3539(WX10234,WX9656,WX10235);
  and AND2_3540(WX10240,WX10239,WX10056);
  and AND2_3541(WX10241,WX9657,WX10242);
  and AND2_3542(WX10247,WX10246,WX10056);
  and AND2_3543(WX10248,WX9658,WX10249);
  and AND2_3544(WX10254,WX10253,WX10056);
  and AND2_3545(WX10255,WX9659,WX10256);
  and AND2_3546(WX10261,WX10260,WX10056);
  and AND2_3547(WX10262,WX9660,WX10263);
  and AND2_3548(WX10268,WX10267,WX10056);
  and AND2_3549(WX10269,WX9661,WX10270);
  and AND2_3550(WX10275,WX10274,WX10056);
  and AND2_3551(WX10276,WX9662,WX10277);
  and AND2_3552(WX10315,WX10285,WX10314);
  and AND2_3553(WX10317,WX10313,WX10314);
  and AND2_3554(WX10319,WX10312,WX10314);
  and AND2_3555(WX10321,WX10311,WX10314);
  and AND2_3556(WX10323,WX10284,WX10314);
  and AND2_3557(WX10325,WX10310,WX10314);
  and AND2_3558(WX10327,WX10309,WX10314);
  and AND2_3559(WX10329,WX10308,WX10314);
  and AND2_3560(WX10331,WX10307,WX10314);
  and AND2_3561(WX10333,WX10306,WX10314);
  and AND2_3562(WX10335,WX10305,WX10314);
  and AND2_3563(WX10337,WX10283,WX10314);
  and AND2_3564(WX10339,WX10304,WX10314);
  and AND2_3565(WX10341,WX10303,WX10314);
  and AND2_3566(WX10343,WX10302,WX10314);
  and AND2_3567(WX10345,WX10301,WX10314);
  and AND2_3568(WX10347,WX10282,WX10314);
  and AND2_3569(WX10349,WX10300,WX10314);
  and AND2_3570(WX10351,WX10299,WX10314);
  and AND2_3571(WX10353,WX10298,WX10314);
  and AND2_3572(WX10355,WX10297,WX10314);
  and AND2_3573(WX10357,WX10296,WX10314);
  and AND2_3574(WX10359,WX10295,WX10314);
  and AND2_3575(WX10361,WX10294,WX10314);
  and AND2_3576(WX10363,WX10293,WX10314);
  and AND2_3577(WX10365,WX10292,WX10314);
  and AND2_3578(WX10367,WX10291,WX10314);
  and AND2_3579(WX10369,WX10290,WX10314);
  and AND2_3580(WX10371,WX10289,WX10314);
  and AND2_3581(WX10373,WX10288,WX10314);
  and AND2_3582(WX10375,WX10287,WX10314);
  and AND2_3583(WX10377,WX10286,WX10314);
  and AND2_3584(WX10379,WX10390,WX11347);
  and AND2_3585(WX10380,WX10386,WX10381);
  and AND2_3586(WX10383,CRC_OUT_1_31,WX11348);
  and AND2_3587(WX10384,DATA_0_31,WX10385);
  and AND2_3588(WX10387,WX10829,WX11348);
  and AND2_3589(WX10388,WX11356,WX10389);
  and AND2_3590(WX10393,WX10404,WX11347);
  and AND2_3591(WX10394,WX10400,WX10395);
  and AND2_3592(WX10397,CRC_OUT_1_30,WX11348);
  and AND2_3593(WX10398,DATA_0_30,WX10399);
  and AND2_3594(WX10401,WX10831,WX11348);
  and AND2_3595(WX10402,WX11363,WX10403);
  and AND2_3596(WX10407,WX10418,WX11347);
  and AND2_3597(WX10408,WX10414,WX10409);
  and AND2_3598(WX10411,CRC_OUT_1_29,WX11348);
  and AND2_3599(WX10412,DATA_0_29,WX10413);
  and AND2_3600(WX10415,WX10833,WX11348);
  and AND2_3601(WX10416,WX11370,WX10417);
  and AND2_3602(WX10421,WX10432,WX11347);
  and AND2_3603(WX10422,WX10428,WX10423);
  and AND2_3604(WX10425,CRC_OUT_1_28,WX11348);
  and AND2_3605(WX10426,DATA_0_28,WX10427);
  and AND2_3606(WX10429,WX10835,WX11348);
  and AND2_3607(WX10430,WX11377,WX10431);
  and AND2_3608(WX10435,WX10446,WX11347);
  and AND2_3609(WX10436,WX10442,WX10437);
  and AND2_3610(WX10439,CRC_OUT_1_27,WX11348);
  and AND2_3611(WX10440,DATA_0_27,WX10441);
  and AND2_3612(WX10443,WX10837,WX11348);
  and AND2_3613(WX10444,WX11384,WX10445);
  and AND2_3614(WX10449,WX10460,WX11347);
  and AND2_3615(WX10450,WX10456,WX10451);
  and AND2_3616(WX10453,CRC_OUT_1_26,WX11348);
  and AND2_3617(WX10454,DATA_0_26,WX10455);
  and AND2_3618(WX10457,WX10839,WX11348);
  and AND2_3619(WX10458,WX11391,WX10459);
  and AND2_3620(WX10463,WX10474,WX11347);
  and AND2_3621(WX10464,WX10470,WX10465);
  and AND2_3622(WX10467,CRC_OUT_1_25,WX11348);
  and AND2_3623(WX10468,DATA_0_25,WX10469);
  and AND2_3624(WX10471,WX10841,WX11348);
  and AND2_3625(WX10472,WX11398,WX10473);
  and AND2_3626(WX10477,WX10488,WX11347);
  and AND2_3627(WX10478,WX10484,WX10479);
  and AND2_3628(WX10481,CRC_OUT_1_24,WX11348);
  and AND2_3629(WX10482,DATA_0_24,WX10483);
  and AND2_3630(WX10485,WX10843,WX11348);
  and AND2_3631(WX10486,WX11405,WX10487);
  and AND2_3632(WX10491,WX10502,WX11347);
  and AND2_3633(WX10492,WX10498,WX10493);
  and AND2_3634(WX10495,CRC_OUT_1_23,WX11348);
  and AND2_3635(WX10496,DATA_0_23,WX10497);
  and AND2_3636(WX10499,WX10845,WX11348);
  and AND2_3637(WX10500,WX11412,WX10501);
  and AND2_3638(WX10505,WX10516,WX11347);
  and AND2_3639(WX10506,WX10512,WX10507);
  and AND2_3640(WX10509,CRC_OUT_1_22,WX11348);
  and AND2_3641(WX10510,DATA_0_22,WX10511);
  and AND2_3642(WX10513,WX10847,WX11348);
  and AND2_3643(WX10514,WX11419,WX10515);
  and AND2_3644(WX10519,WX10530,WX11347);
  and AND2_3645(WX10520,WX10526,WX10521);
  and AND2_3646(WX10523,CRC_OUT_1_21,WX11348);
  and AND2_3647(WX10524,DATA_0_21,WX10525);
  and AND2_3648(WX10527,WX10849,WX11348);
  and AND2_3649(WX10528,WX11426,WX10529);
  and AND2_3650(WX10533,WX10544,WX11347);
  and AND2_3651(WX10534,WX10540,WX10535);
  and AND2_3652(WX10537,CRC_OUT_1_20,WX11348);
  and AND2_3653(WX10538,DATA_0_20,WX10539);
  and AND2_3654(WX10541,WX10851,WX11348);
  and AND2_3655(WX10542,WX11433,WX10543);
  and AND2_3656(WX10547,WX10558,WX11347);
  and AND2_3657(WX10548,WX10554,WX10549);
  and AND2_3658(WX10551,CRC_OUT_1_19,WX11348);
  and AND2_3659(WX10552,DATA_0_19,WX10553);
  and AND2_3660(WX10555,WX10853,WX11348);
  and AND2_3661(WX10556,WX11440,WX10557);
  and AND2_3662(WX10561,WX10572,WX11347);
  and AND2_3663(WX10562,WX10568,WX10563);
  and AND2_3664(WX10565,CRC_OUT_1_18,WX11348);
  and AND2_3665(WX10566,DATA_0_18,WX10567);
  and AND2_3666(WX10569,WX10855,WX11348);
  and AND2_3667(WX10570,WX11447,WX10571);
  and AND2_3668(WX10575,WX10586,WX11347);
  and AND2_3669(WX10576,WX10582,WX10577);
  and AND2_3670(WX10579,CRC_OUT_1_17,WX11348);
  and AND2_3671(WX10580,DATA_0_17,WX10581);
  and AND2_3672(WX10583,WX10857,WX11348);
  and AND2_3673(WX10584,WX11454,WX10585);
  and AND2_3674(WX10589,WX10600,WX11347);
  and AND2_3675(WX10590,WX10596,WX10591);
  and AND2_3676(WX10593,CRC_OUT_1_16,WX11348);
  and AND2_3677(WX10594,DATA_0_16,WX10595);
  and AND2_3678(WX10597,WX10859,WX11348);
  and AND2_3679(WX10598,WX11461,WX10599);
  and AND2_3680(WX10603,WX10614,WX11347);
  and AND2_3681(WX10604,WX10610,WX10605);
  and AND2_3682(WX10607,CRC_OUT_1_15,WX11348);
  and AND2_3683(WX10608,DATA_0_15,WX10609);
  and AND2_3684(WX10611,WX10861,WX11348);
  and AND2_3685(WX10612,WX11468,WX10613);
  and AND2_3686(WX10617,WX10628,WX11347);
  and AND2_3687(WX10618,WX10624,WX10619);
  and AND2_3688(WX10621,CRC_OUT_1_14,WX11348);
  and AND2_3689(WX10622,DATA_0_14,WX10623);
  and AND2_3690(WX10625,WX10863,WX11348);
  and AND2_3691(WX10626,WX11475,WX10627);
  and AND2_3692(WX10631,WX10642,WX11347);
  and AND2_3693(WX10632,WX10638,WX10633);
  and AND2_3694(WX10635,CRC_OUT_1_13,WX11348);
  and AND2_3695(WX10636,DATA_0_13,WX10637);
  and AND2_3696(WX10639,WX10865,WX11348);
  and AND2_3697(WX10640,WX11482,WX10641);
  and AND2_3698(WX10645,WX10656,WX11347);
  and AND2_3699(WX10646,WX10652,WX10647);
  and AND2_3700(WX10649,CRC_OUT_1_12,WX11348);
  and AND2_3701(WX10650,DATA_0_12,WX10651);
  and AND2_3702(WX10653,WX10867,WX11348);
  and AND2_3703(WX10654,WX11489,WX10655);
  and AND2_3704(WX10659,WX10670,WX11347);
  and AND2_3705(WX10660,WX10666,WX10661);
  and AND2_3706(WX10663,CRC_OUT_1_11,WX11348);
  and AND2_3707(WX10664,DATA_0_11,WX10665);
  and AND2_3708(WX10667,WX10869,WX11348);
  and AND2_3709(WX10668,WX11496,WX10669);
  and AND2_3710(WX10673,WX10684,WX11347);
  and AND2_3711(WX10674,WX10680,WX10675);
  and AND2_3712(WX10677,CRC_OUT_1_10,WX11348);
  and AND2_3713(WX10678,DATA_0_10,WX10679);
  and AND2_3714(WX10681,WX10871,WX11348);
  and AND2_3715(WX10682,WX11503,WX10683);
  and AND2_3716(WX10687,WX10698,WX11347);
  and AND2_3717(WX10688,WX10694,WX10689);
  and AND2_3718(WX10691,CRC_OUT_1_9,WX11348);
  and AND2_3719(WX10692,DATA_0_9,WX10693);
  and AND2_3720(WX10695,WX10873,WX11348);
  and AND2_3721(WX10696,WX11510,WX10697);
  and AND2_3722(WX10701,WX10712,WX11347);
  and AND2_3723(WX10702,WX10708,WX10703);
  and AND2_3724(WX10705,CRC_OUT_1_8,WX11348);
  and AND2_3725(WX10706,DATA_0_8,WX10707);
  and AND2_3726(WX10709,WX10875,WX11348);
  and AND2_3727(WX10710,WX11517,WX10711);
  and AND2_3728(WX10715,WX10726,WX11347);
  and AND2_3729(WX10716,WX10722,WX10717);
  and AND2_3730(WX10719,CRC_OUT_1_7,WX11348);
  and AND2_3731(WX10720,DATA_0_7,WX10721);
  and AND2_3732(WX10723,WX10877,WX11348);
  and AND2_3733(WX10724,WX11524,WX10725);
  and AND2_3734(WX10729,WX10740,WX11347);
  and AND2_3735(WX10730,WX10736,WX10731);
  and AND2_3736(WX10733,CRC_OUT_1_6,WX11348);
  and AND2_3737(WX10734,DATA_0_6,WX10735);
  and AND2_3738(WX10737,WX10879,WX11348);
  and AND2_3739(WX10738,WX11531,WX10739);
  and AND2_3740(WX10743,WX10754,WX11347);
  and AND2_3741(WX10744,WX10750,WX10745);
  and AND2_3742(WX10747,CRC_OUT_1_5,WX11348);
  and AND2_3743(WX10748,DATA_0_5,WX10749);
  and AND2_3744(WX10751,WX10881,WX11348);
  and AND2_3745(WX10752,WX11538,WX10753);
  and AND2_3746(WX10757,WX10768,WX11347);
  and AND2_3747(WX10758,WX10764,WX10759);
  and AND2_3748(WX10761,CRC_OUT_1_4,WX11348);
  and AND2_3749(WX10762,DATA_0_4,WX10763);
  and AND2_3750(WX10765,WX10883,WX11348);
  and AND2_3751(WX10766,WX11545,WX10767);
  and AND2_3752(WX10771,WX10782,WX11347);
  and AND2_3753(WX10772,WX10778,WX10773);
  and AND2_3754(WX10775,CRC_OUT_1_3,WX11348);
  and AND2_3755(WX10776,DATA_0_3,WX10777);
  and AND2_3756(WX10779,WX10885,WX11348);
  and AND2_3757(WX10780,WX11552,WX10781);
  and AND2_3758(WX10785,WX10796,WX11347);
  and AND2_3759(WX10786,WX10792,WX10787);
  and AND2_3760(WX10789,CRC_OUT_1_2,WX11348);
  and AND2_3761(WX10790,DATA_0_2,WX10791);
  and AND2_3762(WX10793,WX10887,WX11348);
  and AND2_3763(WX10794,WX11559,WX10795);
  and AND2_3764(WX10799,WX10810,WX11347);
  and AND2_3765(WX10800,WX10806,WX10801);
  and AND2_3766(WX10803,CRC_OUT_1_1,WX11348);
  and AND2_3767(WX10804,DATA_0_1,WX10805);
  and AND2_3768(WX10807,WX10889,WX11348);
  and AND2_3769(WX10808,WX11566,WX10809);
  and AND2_3770(WX10813,WX10824,WX11347);
  and AND2_3771(WX10814,WX10820,WX10815);
  and AND2_3772(WX10817,CRC_OUT_1_0,WX11348);
  and AND2_3773(WX10818,DATA_0_0,WX10819);
  and AND2_3774(WX10821,WX10891,WX11348);
  and AND2_3775(WX10822,WX11573,WX10823);
  and AND2_3776(WX10828,WX10831,RESET);
  and AND2_3777(WX10830,WX10833,RESET);
  and AND2_3778(WX10832,WX10835,RESET);
  and AND2_3779(WX10834,WX10837,RESET);
  and AND2_3780(WX10836,WX10839,RESET);
  and AND2_3781(WX10838,WX10841,RESET);
  and AND2_3782(WX10840,WX10843,RESET);
  and AND2_3783(WX10842,WX10845,RESET);
  and AND2_3784(WX10844,WX10847,RESET);
  and AND2_3785(WX10846,WX10849,RESET);
  and AND2_3786(WX10848,WX10851,RESET);
  and AND2_3787(WX10850,WX10853,RESET);
  and AND2_3788(WX10852,WX10855,RESET);
  and AND2_3789(WX10854,WX10857,RESET);
  and AND2_3790(WX10856,WX10859,RESET);
  and AND2_3791(WX10858,WX10861,RESET);
  and AND2_3792(WX10860,WX10863,RESET);
  and AND2_3793(WX10862,WX10865,RESET);
  and AND2_3794(WX10864,WX10867,RESET);
  and AND2_3795(WX10866,WX10869,RESET);
  and AND2_3796(WX10868,WX10871,RESET);
  and AND2_3797(WX10870,WX10873,RESET);
  and AND2_3798(WX10872,WX10875,RESET);
  and AND2_3799(WX10874,WX10877,RESET);
  and AND2_3800(WX10876,WX10879,RESET);
  and AND2_3801(WX10878,WX10881,RESET);
  and AND2_3802(WX10880,WX10883,RESET);
  and AND2_3803(WX10882,WX10885,RESET);
  and AND2_3804(WX10884,WX10887,RESET);
  and AND2_3805(WX10886,WX10889,RESET);
  and AND2_3806(WX10888,WX10891,RESET);
  and AND2_3807(WX10890,WX10827,RESET);
  and AND2_3808(WX10988,WX10392,RESET);
  and AND2_3809(WX10990,WX10406,RESET);
  and AND2_3810(WX10992,WX10420,RESET);
  and AND2_3811(WX10994,WX10434,RESET);
  and AND2_3812(WX10996,WX10448,RESET);
  and AND2_3813(WX10998,WX10462,RESET);
  and AND2_3814(WX11000,WX10476,RESET);
  and AND2_3815(WX11002,WX10490,RESET);
  and AND2_3816(WX11004,WX10504,RESET);
  and AND2_3817(WX11006,WX10518,RESET);
  and AND2_3818(WX11008,WX10532,RESET);
  and AND2_3819(WX11010,WX10546,RESET);
  and AND2_3820(WX11012,WX10560,RESET);
  and AND2_3821(WX11014,WX10574,RESET);
  and AND2_3822(WX11016,WX10588,RESET);
  and AND2_3823(WX11018,WX10602,RESET);
  and AND2_3824(WX11020,WX10616,RESET);
  and AND2_3825(WX11022,WX10630,RESET);
  and AND2_3826(WX11024,WX10644,RESET);
  and AND2_3827(WX11026,WX10658,RESET);
  and AND2_3828(WX11028,WX10672,RESET);
  and AND2_3829(WX11030,WX10686,RESET);
  and AND2_3830(WX11032,WX10700,RESET);
  and AND2_3831(WX11034,WX10714,RESET);
  and AND2_3832(WX11036,WX10728,RESET);
  and AND2_3833(WX11038,WX10742,RESET);
  and AND2_3834(WX11040,WX10756,RESET);
  and AND2_3835(WX11042,WX10770,RESET);
  and AND2_3836(WX11044,WX10784,RESET);
  and AND2_3837(WX11046,WX10798,RESET);
  and AND2_3838(WX11048,WX10812,RESET);
  and AND2_3839(WX11050,WX10826,RESET);
  and AND2_3840(WX11052,WX10989,RESET);
  and AND2_3841(WX11054,WX10991,RESET);
  and AND2_3842(WX11056,WX10993,RESET);
  and AND2_3843(WX11058,WX10995,RESET);
  and AND2_3844(WX11060,WX10997,RESET);
  and AND2_3845(WX11062,WX10999,RESET);
  and AND2_3846(WX11064,WX11001,RESET);
  and AND2_3847(WX11066,WX11003,RESET);
  and AND2_3848(WX11068,WX11005,RESET);
  and AND2_3849(WX11070,WX11007,RESET);
  and AND2_3850(WX11072,WX11009,RESET);
  and AND2_3851(WX11074,WX11011,RESET);
  and AND2_3852(WX11076,WX11013,RESET);
  and AND2_3853(WX11078,WX11015,RESET);
  and AND2_3854(WX11080,WX11017,RESET);
  and AND2_3855(WX11082,WX11019,RESET);
  and AND2_3856(WX11084,WX11021,RESET);
  and AND2_3857(WX11086,WX11023,RESET);
  and AND2_3858(WX11088,WX11025,RESET);
  and AND2_3859(WX11090,WX11027,RESET);
  and AND2_3860(WX11092,WX11029,RESET);
  and AND2_3861(WX11094,WX11031,RESET);
  and AND2_3862(WX11096,WX11033,RESET);
  and AND2_3863(WX11098,WX11035,RESET);
  and AND2_3864(WX11100,WX11037,RESET);
  and AND2_3865(WX11102,WX11039,RESET);
  and AND2_3866(WX11104,WX11041,RESET);
  and AND2_3867(WX11106,WX11043,RESET);
  and AND2_3868(WX11108,WX11045,RESET);
  and AND2_3869(WX11110,WX11047,RESET);
  and AND2_3870(WX11112,WX11049,RESET);
  and AND2_3871(WX11114,WX11051,RESET);
  and AND2_3872(WX11116,WX11053,RESET);
  and AND2_3873(WX11118,WX11055,RESET);
  and AND2_3874(WX11120,WX11057,RESET);
  and AND2_3875(WX11122,WX11059,RESET);
  and AND2_3876(WX11124,WX11061,RESET);
  and AND2_3877(WX11126,WX11063,RESET);
  and AND2_3878(WX11128,WX11065,RESET);
  and AND2_3879(WX11130,WX11067,RESET);
  and AND2_3880(WX11132,WX11069,RESET);
  and AND2_3881(WX11134,WX11071,RESET);
  and AND2_3882(WX11136,WX11073,RESET);
  and AND2_3883(WX11138,WX11075,RESET);
  and AND2_3884(WX11140,WX11077,RESET);
  and AND2_3885(WX11142,WX11079,RESET);
  and AND2_3886(WX11144,WX11081,RESET);
  and AND2_3887(WX11146,WX11083,RESET);
  and AND2_3888(WX11148,WX11085,RESET);
  and AND2_3889(WX11150,WX11087,RESET);
  and AND2_3890(WX11152,WX11089,RESET);
  and AND2_3891(WX11154,WX11091,RESET);
  and AND2_3892(WX11156,WX11093,RESET);
  and AND2_3893(WX11158,WX11095,RESET);
  and AND2_3894(WX11160,WX11097,RESET);
  and AND2_3895(WX11162,WX11099,RESET);
  and AND2_3896(WX11164,WX11101,RESET);
  and AND2_3897(WX11166,WX11103,RESET);
  and AND2_3898(WX11168,WX11105,RESET);
  and AND2_3899(WX11170,WX11107,RESET);
  and AND2_3900(WX11172,WX11109,RESET);
  and AND2_3901(WX11174,WX11111,RESET);
  and AND2_3902(WX11176,WX11113,RESET);
  and AND2_3903(WX11178,WX11115,RESET);
  and AND2_3904(WX11180,WX11117,RESET);
  and AND2_3905(WX11182,WX11119,RESET);
  and AND2_3906(WX11184,WX11121,RESET);
  and AND2_3907(WX11186,WX11123,RESET);
  and AND2_3908(WX11188,WX11125,RESET);
  and AND2_3909(WX11190,WX11127,RESET);
  and AND2_3910(WX11192,WX11129,RESET);
  and AND2_3911(WX11194,WX11131,RESET);
  and AND2_3912(WX11196,WX11133,RESET);
  and AND2_3913(WX11198,WX11135,RESET);
  and AND2_3914(WX11200,WX11137,RESET);
  and AND2_3915(WX11202,WX11139,RESET);
  and AND2_3916(WX11204,WX11141,RESET);
  and AND2_3917(WX11206,WX11143,RESET);
  and AND2_3918(WX11208,WX11145,RESET);
  and AND2_3919(WX11210,WX11147,RESET);
  and AND2_3920(WX11212,WX11149,RESET);
  and AND2_3921(WX11214,WX11151,RESET);
  and AND2_3922(WX11216,WX11153,RESET);
  and AND2_3923(WX11218,WX11155,RESET);
  and AND2_3924(WX11220,WX11157,RESET);
  and AND2_3925(WX11222,WX11159,RESET);
  and AND2_3926(WX11224,WX11161,RESET);
  and AND2_3927(WX11226,WX11163,RESET);
  and AND2_3928(WX11228,WX11165,RESET);
  and AND2_3929(WX11230,WX11167,RESET);
  and AND2_3930(WX11232,WX11169,RESET);
  and AND2_3931(WX11234,WX11171,RESET);
  and AND2_3932(WX11236,WX11173,RESET);
  and AND2_3933(WX11238,WX11175,RESET);
  and AND2_3934(WX11240,WX11177,RESET);
  and AND2_3935(WX11242,WX11179,RESET);
  and AND2_3936(WX11351,WX11350,WX11349);
  and AND2_3937(WX11352,WX10924,WX11353);
  and AND2_3938(WX11358,WX11357,WX11349);
  and AND2_3939(WX11359,WX10925,WX11360);
  and AND2_3940(WX11365,WX11364,WX11349);
  and AND2_3941(WX11366,WX10926,WX11367);
  and AND2_3942(WX11372,WX11371,WX11349);
  and AND2_3943(WX11373,WX10927,WX11374);
  and AND2_3944(WX11379,WX11378,WX11349);
  and AND2_3945(WX11380,WX10928,WX11381);
  and AND2_3946(WX11386,WX11385,WX11349);
  and AND2_3947(WX11387,WX10929,WX11388);
  and AND2_3948(WX11393,WX11392,WX11349);
  and AND2_3949(WX11394,WX10930,WX11395);
  and AND2_3950(WX11400,WX11399,WX11349);
  and AND2_3951(WX11401,WX10931,WX11402);
  and AND2_3952(WX11407,WX11406,WX11349);
  and AND2_3953(WX11408,WX10932,WX11409);
  and AND2_3954(WX11414,WX11413,WX11349);
  and AND2_3955(WX11415,WX10933,WX11416);
  and AND2_3956(WX11421,WX11420,WX11349);
  and AND2_3957(WX11422,WX10934,WX11423);
  and AND2_3958(WX11428,WX11427,WX11349);
  and AND2_3959(WX11429,WX10935,WX11430);
  and AND2_3960(WX11435,WX11434,WX11349);
  and AND2_3961(WX11436,WX10936,WX11437);
  and AND2_3962(WX11442,WX11441,WX11349);
  and AND2_3963(WX11443,WX10937,WX11444);
  and AND2_3964(WX11449,WX11448,WX11349);
  and AND2_3965(WX11450,WX10938,WX11451);
  and AND2_3966(WX11456,WX11455,WX11349);
  and AND2_3967(WX11457,WX10939,WX11458);
  and AND2_3968(WX11463,WX11462,WX11349);
  and AND2_3969(WX11464,WX10940,WX11465);
  and AND2_3970(WX11470,WX11469,WX11349);
  and AND2_3971(WX11471,WX10941,WX11472);
  and AND2_3972(WX11477,WX11476,WX11349);
  and AND2_3973(WX11478,WX10942,WX11479);
  and AND2_3974(WX11484,WX11483,WX11349);
  and AND2_3975(WX11485,WX10943,WX11486);
  and AND2_3976(WX11491,WX11490,WX11349);
  and AND2_3977(WX11492,WX10944,WX11493);
  and AND2_3978(WX11498,WX11497,WX11349);
  and AND2_3979(WX11499,WX10945,WX11500);
  and AND2_3980(WX11505,WX11504,WX11349);
  and AND2_3981(WX11506,WX10946,WX11507);
  and AND2_3982(WX11512,WX11511,WX11349);
  and AND2_3983(WX11513,WX10947,WX11514);
  and AND2_3984(WX11519,WX11518,WX11349);
  and AND2_3985(WX11520,WX10948,WX11521);
  and AND2_3986(WX11526,WX11525,WX11349);
  and AND2_3987(WX11527,WX10949,WX11528);
  and AND2_3988(WX11533,WX11532,WX11349);
  and AND2_3989(WX11534,WX10950,WX11535);
  and AND2_3990(WX11540,WX11539,WX11349);
  and AND2_3991(WX11541,WX10951,WX11542);
  and AND2_3992(WX11547,WX11546,WX11349);
  and AND2_3993(WX11548,WX10952,WX11549);
  and AND2_3994(WX11554,WX11553,WX11349);
  and AND2_3995(WX11555,WX10953,WX11556);
  and AND2_3996(WX11561,WX11560,WX11349);
  and AND2_3997(WX11562,WX10954,WX11563);
  and AND2_3998(WX11568,WX11567,WX11349);
  and AND2_3999(WX11569,WX10955,WX11570);
  and AND2_4000(WX11608,WX11578,WX11607);
  and AND2_4001(WX11610,WX11606,WX11607);
  and AND2_4002(WX11612,WX11605,WX11607);
  and AND2_4003(WX11614,WX11604,WX11607);
  and AND2_4004(WX11616,WX11577,WX11607);
  and AND2_4005(WX11618,WX11603,WX11607);
  and AND2_4006(WX11620,WX11602,WX11607);
  and AND2_4007(WX11622,WX11601,WX11607);
  and AND2_4008(WX11624,WX11600,WX11607);
  and AND2_4009(WX11626,WX11599,WX11607);
  and AND2_4010(WX11628,WX11598,WX11607);
  and AND2_4011(WX11630,WX11576,WX11607);
  and AND2_4012(WX11632,WX11597,WX11607);
  and AND2_4013(WX11634,WX11596,WX11607);
  and AND2_4014(WX11636,WX11595,WX11607);
  and AND2_4015(WX11638,WX11594,WX11607);
  and AND2_4016(WX11640,WX11575,WX11607);
  and AND2_4017(WX11642,WX11593,WX11607);
  and AND2_4018(WX11644,WX11592,WX11607);
  and AND2_4019(WX11646,WX11591,WX11607);
  and AND2_4020(WX11648,WX11590,WX11607);
  and AND2_4021(WX11650,WX11589,WX11607);
  and AND2_4022(WX11652,WX11588,WX11607);
  and AND2_4023(WX11654,WX11587,WX11607);
  and AND2_4024(WX11656,WX11586,WX11607);
  and AND2_4025(WX11658,WX11585,WX11607);
  and AND2_4026(WX11660,WX11584,WX11607);
  and AND2_4027(WX11662,WX11583,WX11607);
  and AND2_4028(WX11664,WX11582,WX11607);
  and AND2_4029(WX11666,WX11581,WX11607);
  and AND2_4030(WX11668,WX11580,WX11607);
  and AND2_4031(WX11670,WX11579,WX11607);
  or OR2_0(WX38,WX36,WX35);
  or OR2_1(WX42,WX40,WX39);
  or OR2_2(WX46,WX44,WX43);
  or OR2_3(WX52,WX50,WX49);
  or OR2_4(WX56,WX54,WX53);
  or OR2_5(WX60,WX58,WX57);
  or OR2_6(WX66,WX64,WX63);
  or OR2_7(WX70,WX68,WX67);
  or OR2_8(WX74,WX72,WX71);
  or OR2_9(WX80,WX78,WX77);
  or OR2_10(WX84,WX82,WX81);
  or OR2_11(WX88,WX86,WX85);
  or OR2_12(WX94,WX92,WX91);
  or OR2_13(WX98,WX96,WX95);
  or OR2_14(WX102,WX100,WX99);
  or OR2_15(WX108,WX106,WX105);
  or OR2_16(WX112,WX110,WX109);
  or OR2_17(WX116,WX114,WX113);
  or OR2_18(WX122,WX120,WX119);
  or OR2_19(WX126,WX124,WX123);
  or OR2_20(WX130,WX128,WX127);
  or OR2_21(WX136,WX134,WX133);
  or OR2_22(WX140,WX138,WX137);
  or OR2_23(WX144,WX142,WX141);
  or OR2_24(WX150,WX148,WX147);
  or OR2_25(WX154,WX152,WX151);
  or OR2_26(WX158,WX156,WX155);
  or OR2_27(WX164,WX162,WX161);
  or OR2_28(WX168,WX166,WX165);
  or OR2_29(WX172,WX170,WX169);
  or OR2_30(WX178,WX176,WX175);
  or OR2_31(WX182,WX180,WX179);
  or OR2_32(WX186,WX184,WX183);
  or OR2_33(WX192,WX190,WX189);
  or OR2_34(WX196,WX194,WX193);
  or OR2_35(WX200,WX198,WX197);
  or OR2_36(WX206,WX204,WX203);
  or OR2_37(WX210,WX208,WX207);
  or OR2_38(WX214,WX212,WX211);
  or OR2_39(WX220,WX218,WX217);
  or OR2_40(WX224,WX222,WX221);
  or OR2_41(WX228,WX226,WX225);
  or OR2_42(WX234,WX232,WX231);
  or OR2_43(WX238,WX236,WX235);
  or OR2_44(WX242,WX240,WX239);
  or OR2_45(WX248,WX246,WX245);
  or OR2_46(WX252,WX250,WX249);
  or OR2_47(WX256,WX254,WX253);
  or OR2_48(WX262,WX260,WX259);
  or OR2_49(WX266,WX264,WX263);
  or OR2_50(WX270,WX268,WX267);
  or OR2_51(WX276,WX274,WX273);
  or OR2_52(WX280,WX278,WX277);
  or OR2_53(WX284,WX282,WX281);
  or OR2_54(WX290,WX288,WX287);
  or OR2_55(WX294,WX292,WX291);
  or OR2_56(WX298,WX296,WX295);
  or OR2_57(WX304,WX302,WX301);
  or OR2_58(WX308,WX306,WX305);
  or OR2_59(WX312,WX310,WX309);
  or OR2_60(WX318,WX316,WX315);
  or OR2_61(WX322,WX320,WX319);
  or OR2_62(WX326,WX324,WX323);
  or OR2_63(WX332,WX330,WX329);
  or OR2_64(WX336,WX334,WX333);
  or OR2_65(WX340,WX338,WX337);
  or OR2_66(WX346,WX344,WX343);
  or OR2_67(WX350,WX348,WX347);
  or OR2_68(WX354,WX352,WX351);
  or OR2_69(WX360,WX358,WX357);
  or OR2_70(WX364,WX362,WX361);
  or OR2_71(WX368,WX366,WX365);
  or OR2_72(WX374,WX372,WX371);
  or OR2_73(WX378,WX376,WX375);
  or OR2_74(WX382,WX380,WX379);
  or OR2_75(WX388,WX386,WX385);
  or OR2_76(WX392,WX390,WX389);
  or OR2_77(WX396,WX394,WX393);
  or OR2_78(WX402,WX400,WX399);
  or OR2_79(WX406,WX404,WX403);
  or OR2_80(WX410,WX408,WX407);
  or OR2_81(WX416,WX414,WX413);
  or OR2_82(WX420,WX418,WX417);
  or OR2_83(WX424,WX422,WX421);
  or OR2_84(WX430,WX428,WX427);
  or OR2_85(WX434,WX432,WX431);
  or OR2_86(WX438,WX436,WX435);
  or OR2_87(WX444,WX442,WX441);
  or OR2_88(WX448,WX446,WX445);
  or OR2_89(WX452,WX450,WX449);
  or OR2_90(WX458,WX456,WX455);
  or OR2_91(WX462,WX460,WX459);
  or OR2_92(WX466,WX464,WX463);
  or OR2_93(WX472,WX470,WX469);
  or OR2_94(WX476,WX474,WX473);
  or OR2_95(WX480,WX478,WX477);
  or OR2_96(WX1010,WX1008,WX1007);
  or OR2_97(WX1017,WX1015,WX1014);
  or OR2_98(WX1024,WX1022,WX1021);
  or OR2_99(WX1031,WX1029,WX1028);
  or OR2_100(WX1038,WX1036,WX1035);
  or OR2_101(WX1045,WX1043,WX1042);
  or OR2_102(WX1052,WX1050,WX1049);
  or OR2_103(WX1059,WX1057,WX1056);
  or OR2_104(WX1066,WX1064,WX1063);
  or OR2_105(WX1073,WX1071,WX1070);
  or OR2_106(WX1080,WX1078,WX1077);
  or OR2_107(WX1087,WX1085,WX1084);
  or OR2_108(WX1094,WX1092,WX1091);
  or OR2_109(WX1101,WX1099,WX1098);
  or OR2_110(WX1108,WX1106,WX1105);
  or OR2_111(WX1115,WX1113,WX1112);
  or OR2_112(WX1122,WX1120,WX1119);
  or OR2_113(WX1129,WX1127,WX1126);
  or OR2_114(WX1136,WX1134,WX1133);
  or OR2_115(WX1143,WX1141,WX1140);
  or OR2_116(WX1150,WX1148,WX1147);
  or OR2_117(WX1157,WX1155,WX1154);
  or OR2_118(WX1164,WX1162,WX1161);
  or OR2_119(WX1171,WX1169,WX1168);
  or OR2_120(WX1178,WX1176,WX1175);
  or OR2_121(WX1185,WX1183,WX1182);
  or OR2_122(WX1192,WX1190,WX1189);
  or OR2_123(WX1199,WX1197,WX1196);
  or OR2_124(WX1206,WX1204,WX1203);
  or OR2_125(WX1213,WX1211,WX1210);
  or OR2_126(WX1220,WX1218,WX1217);
  or OR2_127(WX1227,WX1225,WX1224);
  or OR2_128(WX1331,WX1329,WX1328);
  or OR2_129(WX1335,WX1333,WX1332);
  or OR2_130(WX1339,WX1337,WX1336);
  or OR2_131(WX1345,WX1343,WX1342);
  or OR2_132(WX1349,WX1347,WX1346);
  or OR2_133(WX1353,WX1351,WX1350);
  or OR2_134(WX1359,WX1357,WX1356);
  or OR2_135(WX1363,WX1361,WX1360);
  or OR2_136(WX1367,WX1365,WX1364);
  or OR2_137(WX1373,WX1371,WX1370);
  or OR2_138(WX1377,WX1375,WX1374);
  or OR2_139(WX1381,WX1379,WX1378);
  or OR2_140(WX1387,WX1385,WX1384);
  or OR2_141(WX1391,WX1389,WX1388);
  or OR2_142(WX1395,WX1393,WX1392);
  or OR2_143(WX1401,WX1399,WX1398);
  or OR2_144(WX1405,WX1403,WX1402);
  or OR2_145(WX1409,WX1407,WX1406);
  or OR2_146(WX1415,WX1413,WX1412);
  or OR2_147(WX1419,WX1417,WX1416);
  or OR2_148(WX1423,WX1421,WX1420);
  or OR2_149(WX1429,WX1427,WX1426);
  or OR2_150(WX1433,WX1431,WX1430);
  or OR2_151(WX1437,WX1435,WX1434);
  or OR2_152(WX1443,WX1441,WX1440);
  or OR2_153(WX1447,WX1445,WX1444);
  or OR2_154(WX1451,WX1449,WX1448);
  or OR2_155(WX1457,WX1455,WX1454);
  or OR2_156(WX1461,WX1459,WX1458);
  or OR2_157(WX1465,WX1463,WX1462);
  or OR2_158(WX1471,WX1469,WX1468);
  or OR2_159(WX1475,WX1473,WX1472);
  or OR2_160(WX1479,WX1477,WX1476);
  or OR2_161(WX1485,WX1483,WX1482);
  or OR2_162(WX1489,WX1487,WX1486);
  or OR2_163(WX1493,WX1491,WX1490);
  or OR2_164(WX1499,WX1497,WX1496);
  or OR2_165(WX1503,WX1501,WX1500);
  or OR2_166(WX1507,WX1505,WX1504);
  or OR2_167(WX1513,WX1511,WX1510);
  or OR2_168(WX1517,WX1515,WX1514);
  or OR2_169(WX1521,WX1519,WX1518);
  or OR2_170(WX1527,WX1525,WX1524);
  or OR2_171(WX1531,WX1529,WX1528);
  or OR2_172(WX1535,WX1533,WX1532);
  or OR2_173(WX1541,WX1539,WX1538);
  or OR2_174(WX1545,WX1543,WX1542);
  or OR2_175(WX1549,WX1547,WX1546);
  or OR2_176(WX1555,WX1553,WX1552);
  or OR2_177(WX1559,WX1557,WX1556);
  or OR2_178(WX1563,WX1561,WX1560);
  or OR2_179(WX1569,WX1567,WX1566);
  or OR2_180(WX1573,WX1571,WX1570);
  or OR2_181(WX1577,WX1575,WX1574);
  or OR2_182(WX1583,WX1581,WX1580);
  or OR2_183(WX1587,WX1585,WX1584);
  or OR2_184(WX1591,WX1589,WX1588);
  or OR2_185(WX1597,WX1595,WX1594);
  or OR2_186(WX1601,WX1599,WX1598);
  or OR2_187(WX1605,WX1603,WX1602);
  or OR2_188(WX1611,WX1609,WX1608);
  or OR2_189(WX1615,WX1613,WX1612);
  or OR2_190(WX1619,WX1617,WX1616);
  or OR2_191(WX1625,WX1623,WX1622);
  or OR2_192(WX1629,WX1627,WX1626);
  or OR2_193(WX1633,WX1631,WX1630);
  or OR2_194(WX1639,WX1637,WX1636);
  or OR2_195(WX1643,WX1641,WX1640);
  or OR2_196(WX1647,WX1645,WX1644);
  or OR2_197(WX1653,WX1651,WX1650);
  or OR2_198(WX1657,WX1655,WX1654);
  or OR2_199(WX1661,WX1659,WX1658);
  or OR2_200(WX1667,WX1665,WX1664);
  or OR2_201(WX1671,WX1669,WX1668);
  or OR2_202(WX1675,WX1673,WX1672);
  or OR2_203(WX1681,WX1679,WX1678);
  or OR2_204(WX1685,WX1683,WX1682);
  or OR2_205(WX1689,WX1687,WX1686);
  or OR2_206(WX1695,WX1693,WX1692);
  or OR2_207(WX1699,WX1697,WX1696);
  or OR2_208(WX1703,WX1701,WX1700);
  or OR2_209(WX1709,WX1707,WX1706);
  or OR2_210(WX1713,WX1711,WX1710);
  or OR2_211(WX1717,WX1715,WX1714);
  or OR2_212(WX1723,WX1721,WX1720);
  or OR2_213(WX1727,WX1725,WX1724);
  or OR2_214(WX1731,WX1729,WX1728);
  or OR2_215(WX1737,WX1735,WX1734);
  or OR2_216(WX1741,WX1739,WX1738);
  or OR2_217(WX1745,WX1743,WX1742);
  or OR2_218(WX1751,WX1749,WX1748);
  or OR2_219(WX1755,WX1753,WX1752);
  or OR2_220(WX1759,WX1757,WX1756);
  or OR2_221(WX1765,WX1763,WX1762);
  or OR2_222(WX1769,WX1767,WX1766);
  or OR2_223(WX1773,WX1771,WX1770);
  or OR2_224(WX2303,WX2301,WX2300);
  or OR2_225(WX2310,WX2308,WX2307);
  or OR2_226(WX2317,WX2315,WX2314);
  or OR2_227(WX2324,WX2322,WX2321);
  or OR2_228(WX2331,WX2329,WX2328);
  or OR2_229(WX2338,WX2336,WX2335);
  or OR2_230(WX2345,WX2343,WX2342);
  or OR2_231(WX2352,WX2350,WX2349);
  or OR2_232(WX2359,WX2357,WX2356);
  or OR2_233(WX2366,WX2364,WX2363);
  or OR2_234(WX2373,WX2371,WX2370);
  or OR2_235(WX2380,WX2378,WX2377);
  or OR2_236(WX2387,WX2385,WX2384);
  or OR2_237(WX2394,WX2392,WX2391);
  or OR2_238(WX2401,WX2399,WX2398);
  or OR2_239(WX2408,WX2406,WX2405);
  or OR2_240(WX2415,WX2413,WX2412);
  or OR2_241(WX2422,WX2420,WX2419);
  or OR2_242(WX2429,WX2427,WX2426);
  or OR2_243(WX2436,WX2434,WX2433);
  or OR2_244(WX2443,WX2441,WX2440);
  or OR2_245(WX2450,WX2448,WX2447);
  or OR2_246(WX2457,WX2455,WX2454);
  or OR2_247(WX2464,WX2462,WX2461);
  or OR2_248(WX2471,WX2469,WX2468);
  or OR2_249(WX2478,WX2476,WX2475);
  or OR2_250(WX2485,WX2483,WX2482);
  or OR2_251(WX2492,WX2490,WX2489);
  or OR2_252(WX2499,WX2497,WX2496);
  or OR2_253(WX2506,WX2504,WX2503);
  or OR2_254(WX2513,WX2511,WX2510);
  or OR2_255(WX2520,WX2518,WX2517);
  or OR2_256(WX2624,WX2622,WX2621);
  or OR2_257(WX2628,WX2626,WX2625);
  or OR2_258(WX2632,WX2630,WX2629);
  or OR2_259(WX2638,WX2636,WX2635);
  or OR2_260(WX2642,WX2640,WX2639);
  or OR2_261(WX2646,WX2644,WX2643);
  or OR2_262(WX2652,WX2650,WX2649);
  or OR2_263(WX2656,WX2654,WX2653);
  or OR2_264(WX2660,WX2658,WX2657);
  or OR2_265(WX2666,WX2664,WX2663);
  or OR2_266(WX2670,WX2668,WX2667);
  or OR2_267(WX2674,WX2672,WX2671);
  or OR2_268(WX2680,WX2678,WX2677);
  or OR2_269(WX2684,WX2682,WX2681);
  or OR2_270(WX2688,WX2686,WX2685);
  or OR2_271(WX2694,WX2692,WX2691);
  or OR2_272(WX2698,WX2696,WX2695);
  or OR2_273(WX2702,WX2700,WX2699);
  or OR2_274(WX2708,WX2706,WX2705);
  or OR2_275(WX2712,WX2710,WX2709);
  or OR2_276(WX2716,WX2714,WX2713);
  or OR2_277(WX2722,WX2720,WX2719);
  or OR2_278(WX2726,WX2724,WX2723);
  or OR2_279(WX2730,WX2728,WX2727);
  or OR2_280(WX2736,WX2734,WX2733);
  or OR2_281(WX2740,WX2738,WX2737);
  or OR2_282(WX2744,WX2742,WX2741);
  or OR2_283(WX2750,WX2748,WX2747);
  or OR2_284(WX2754,WX2752,WX2751);
  or OR2_285(WX2758,WX2756,WX2755);
  or OR2_286(WX2764,WX2762,WX2761);
  or OR2_287(WX2768,WX2766,WX2765);
  or OR2_288(WX2772,WX2770,WX2769);
  or OR2_289(WX2778,WX2776,WX2775);
  or OR2_290(WX2782,WX2780,WX2779);
  or OR2_291(WX2786,WX2784,WX2783);
  or OR2_292(WX2792,WX2790,WX2789);
  or OR2_293(WX2796,WX2794,WX2793);
  or OR2_294(WX2800,WX2798,WX2797);
  or OR2_295(WX2806,WX2804,WX2803);
  or OR2_296(WX2810,WX2808,WX2807);
  or OR2_297(WX2814,WX2812,WX2811);
  or OR2_298(WX2820,WX2818,WX2817);
  or OR2_299(WX2824,WX2822,WX2821);
  or OR2_300(WX2828,WX2826,WX2825);
  or OR2_301(WX2834,WX2832,WX2831);
  or OR2_302(WX2838,WX2836,WX2835);
  or OR2_303(WX2842,WX2840,WX2839);
  or OR2_304(WX2848,WX2846,WX2845);
  or OR2_305(WX2852,WX2850,WX2849);
  or OR2_306(WX2856,WX2854,WX2853);
  or OR2_307(WX2862,WX2860,WX2859);
  or OR2_308(WX2866,WX2864,WX2863);
  or OR2_309(WX2870,WX2868,WX2867);
  or OR2_310(WX2876,WX2874,WX2873);
  or OR2_311(WX2880,WX2878,WX2877);
  or OR2_312(WX2884,WX2882,WX2881);
  or OR2_313(WX2890,WX2888,WX2887);
  or OR2_314(WX2894,WX2892,WX2891);
  or OR2_315(WX2898,WX2896,WX2895);
  or OR2_316(WX2904,WX2902,WX2901);
  or OR2_317(WX2908,WX2906,WX2905);
  or OR2_318(WX2912,WX2910,WX2909);
  or OR2_319(WX2918,WX2916,WX2915);
  or OR2_320(WX2922,WX2920,WX2919);
  or OR2_321(WX2926,WX2924,WX2923);
  or OR2_322(WX2932,WX2930,WX2929);
  or OR2_323(WX2936,WX2934,WX2933);
  or OR2_324(WX2940,WX2938,WX2937);
  or OR2_325(WX2946,WX2944,WX2943);
  or OR2_326(WX2950,WX2948,WX2947);
  or OR2_327(WX2954,WX2952,WX2951);
  or OR2_328(WX2960,WX2958,WX2957);
  or OR2_329(WX2964,WX2962,WX2961);
  or OR2_330(WX2968,WX2966,WX2965);
  or OR2_331(WX2974,WX2972,WX2971);
  or OR2_332(WX2978,WX2976,WX2975);
  or OR2_333(WX2982,WX2980,WX2979);
  or OR2_334(WX2988,WX2986,WX2985);
  or OR2_335(WX2992,WX2990,WX2989);
  or OR2_336(WX2996,WX2994,WX2993);
  or OR2_337(WX3002,WX3000,WX2999);
  or OR2_338(WX3006,WX3004,WX3003);
  or OR2_339(WX3010,WX3008,WX3007);
  or OR2_340(WX3016,WX3014,WX3013);
  or OR2_341(WX3020,WX3018,WX3017);
  or OR2_342(WX3024,WX3022,WX3021);
  or OR2_343(WX3030,WX3028,WX3027);
  or OR2_344(WX3034,WX3032,WX3031);
  or OR2_345(WX3038,WX3036,WX3035);
  or OR2_346(WX3044,WX3042,WX3041);
  or OR2_347(WX3048,WX3046,WX3045);
  or OR2_348(WX3052,WX3050,WX3049);
  or OR2_349(WX3058,WX3056,WX3055);
  or OR2_350(WX3062,WX3060,WX3059);
  or OR2_351(WX3066,WX3064,WX3063);
  or OR2_352(WX3596,WX3594,WX3593);
  or OR2_353(WX3603,WX3601,WX3600);
  or OR2_354(WX3610,WX3608,WX3607);
  or OR2_355(WX3617,WX3615,WX3614);
  or OR2_356(WX3624,WX3622,WX3621);
  or OR2_357(WX3631,WX3629,WX3628);
  or OR2_358(WX3638,WX3636,WX3635);
  or OR2_359(WX3645,WX3643,WX3642);
  or OR2_360(WX3652,WX3650,WX3649);
  or OR2_361(WX3659,WX3657,WX3656);
  or OR2_362(WX3666,WX3664,WX3663);
  or OR2_363(WX3673,WX3671,WX3670);
  or OR2_364(WX3680,WX3678,WX3677);
  or OR2_365(WX3687,WX3685,WX3684);
  or OR2_366(WX3694,WX3692,WX3691);
  or OR2_367(WX3701,WX3699,WX3698);
  or OR2_368(WX3708,WX3706,WX3705);
  or OR2_369(WX3715,WX3713,WX3712);
  or OR2_370(WX3722,WX3720,WX3719);
  or OR2_371(WX3729,WX3727,WX3726);
  or OR2_372(WX3736,WX3734,WX3733);
  or OR2_373(WX3743,WX3741,WX3740);
  or OR2_374(WX3750,WX3748,WX3747);
  or OR2_375(WX3757,WX3755,WX3754);
  or OR2_376(WX3764,WX3762,WX3761);
  or OR2_377(WX3771,WX3769,WX3768);
  or OR2_378(WX3778,WX3776,WX3775);
  or OR2_379(WX3785,WX3783,WX3782);
  or OR2_380(WX3792,WX3790,WX3789);
  or OR2_381(WX3799,WX3797,WX3796);
  or OR2_382(WX3806,WX3804,WX3803);
  or OR2_383(WX3813,WX3811,WX3810);
  or OR2_384(WX3917,WX3915,WX3914);
  or OR2_385(WX3921,WX3919,WX3918);
  or OR2_386(WX3925,WX3923,WX3922);
  or OR2_387(WX3931,WX3929,WX3928);
  or OR2_388(WX3935,WX3933,WX3932);
  or OR2_389(WX3939,WX3937,WX3936);
  or OR2_390(WX3945,WX3943,WX3942);
  or OR2_391(WX3949,WX3947,WX3946);
  or OR2_392(WX3953,WX3951,WX3950);
  or OR2_393(WX3959,WX3957,WX3956);
  or OR2_394(WX3963,WX3961,WX3960);
  or OR2_395(WX3967,WX3965,WX3964);
  or OR2_396(WX3973,WX3971,WX3970);
  or OR2_397(WX3977,WX3975,WX3974);
  or OR2_398(WX3981,WX3979,WX3978);
  or OR2_399(WX3987,WX3985,WX3984);
  or OR2_400(WX3991,WX3989,WX3988);
  or OR2_401(WX3995,WX3993,WX3992);
  or OR2_402(WX4001,WX3999,WX3998);
  or OR2_403(WX4005,WX4003,WX4002);
  or OR2_404(WX4009,WX4007,WX4006);
  or OR2_405(WX4015,WX4013,WX4012);
  or OR2_406(WX4019,WX4017,WX4016);
  or OR2_407(WX4023,WX4021,WX4020);
  or OR2_408(WX4029,WX4027,WX4026);
  or OR2_409(WX4033,WX4031,WX4030);
  or OR2_410(WX4037,WX4035,WX4034);
  or OR2_411(WX4043,WX4041,WX4040);
  or OR2_412(WX4047,WX4045,WX4044);
  or OR2_413(WX4051,WX4049,WX4048);
  or OR2_414(WX4057,WX4055,WX4054);
  or OR2_415(WX4061,WX4059,WX4058);
  or OR2_416(WX4065,WX4063,WX4062);
  or OR2_417(WX4071,WX4069,WX4068);
  or OR2_418(WX4075,WX4073,WX4072);
  or OR2_419(WX4079,WX4077,WX4076);
  or OR2_420(WX4085,WX4083,WX4082);
  or OR2_421(WX4089,WX4087,WX4086);
  or OR2_422(WX4093,WX4091,WX4090);
  or OR2_423(WX4099,WX4097,WX4096);
  or OR2_424(WX4103,WX4101,WX4100);
  or OR2_425(WX4107,WX4105,WX4104);
  or OR2_426(WX4113,WX4111,WX4110);
  or OR2_427(WX4117,WX4115,WX4114);
  or OR2_428(WX4121,WX4119,WX4118);
  or OR2_429(WX4127,WX4125,WX4124);
  or OR2_430(WX4131,WX4129,WX4128);
  or OR2_431(WX4135,WX4133,WX4132);
  or OR2_432(WX4141,WX4139,WX4138);
  or OR2_433(WX4145,WX4143,WX4142);
  or OR2_434(WX4149,WX4147,WX4146);
  or OR2_435(WX4155,WX4153,WX4152);
  or OR2_436(WX4159,WX4157,WX4156);
  or OR2_437(WX4163,WX4161,WX4160);
  or OR2_438(WX4169,WX4167,WX4166);
  or OR2_439(WX4173,WX4171,WX4170);
  or OR2_440(WX4177,WX4175,WX4174);
  or OR2_441(WX4183,WX4181,WX4180);
  or OR2_442(WX4187,WX4185,WX4184);
  or OR2_443(WX4191,WX4189,WX4188);
  or OR2_444(WX4197,WX4195,WX4194);
  or OR2_445(WX4201,WX4199,WX4198);
  or OR2_446(WX4205,WX4203,WX4202);
  or OR2_447(WX4211,WX4209,WX4208);
  or OR2_448(WX4215,WX4213,WX4212);
  or OR2_449(WX4219,WX4217,WX4216);
  or OR2_450(WX4225,WX4223,WX4222);
  or OR2_451(WX4229,WX4227,WX4226);
  or OR2_452(WX4233,WX4231,WX4230);
  or OR2_453(WX4239,WX4237,WX4236);
  or OR2_454(WX4243,WX4241,WX4240);
  or OR2_455(WX4247,WX4245,WX4244);
  or OR2_456(WX4253,WX4251,WX4250);
  or OR2_457(WX4257,WX4255,WX4254);
  or OR2_458(WX4261,WX4259,WX4258);
  or OR2_459(WX4267,WX4265,WX4264);
  or OR2_460(WX4271,WX4269,WX4268);
  or OR2_461(WX4275,WX4273,WX4272);
  or OR2_462(WX4281,WX4279,WX4278);
  or OR2_463(WX4285,WX4283,WX4282);
  or OR2_464(WX4289,WX4287,WX4286);
  or OR2_465(WX4295,WX4293,WX4292);
  or OR2_466(WX4299,WX4297,WX4296);
  or OR2_467(WX4303,WX4301,WX4300);
  or OR2_468(WX4309,WX4307,WX4306);
  or OR2_469(WX4313,WX4311,WX4310);
  or OR2_470(WX4317,WX4315,WX4314);
  or OR2_471(WX4323,WX4321,WX4320);
  or OR2_472(WX4327,WX4325,WX4324);
  or OR2_473(WX4331,WX4329,WX4328);
  or OR2_474(WX4337,WX4335,WX4334);
  or OR2_475(WX4341,WX4339,WX4338);
  or OR2_476(WX4345,WX4343,WX4342);
  or OR2_477(WX4351,WX4349,WX4348);
  or OR2_478(WX4355,WX4353,WX4352);
  or OR2_479(WX4359,WX4357,WX4356);
  or OR2_480(WX4889,WX4887,WX4886);
  or OR2_481(WX4896,WX4894,WX4893);
  or OR2_482(WX4903,WX4901,WX4900);
  or OR2_483(WX4910,WX4908,WX4907);
  or OR2_484(WX4917,WX4915,WX4914);
  or OR2_485(WX4924,WX4922,WX4921);
  or OR2_486(WX4931,WX4929,WX4928);
  or OR2_487(WX4938,WX4936,WX4935);
  or OR2_488(WX4945,WX4943,WX4942);
  or OR2_489(WX4952,WX4950,WX4949);
  or OR2_490(WX4959,WX4957,WX4956);
  or OR2_491(WX4966,WX4964,WX4963);
  or OR2_492(WX4973,WX4971,WX4970);
  or OR2_493(WX4980,WX4978,WX4977);
  or OR2_494(WX4987,WX4985,WX4984);
  or OR2_495(WX4994,WX4992,WX4991);
  or OR2_496(WX5001,WX4999,WX4998);
  or OR2_497(WX5008,WX5006,WX5005);
  or OR2_498(WX5015,WX5013,WX5012);
  or OR2_499(WX5022,WX5020,WX5019);
  or OR2_500(WX5029,WX5027,WX5026);
  or OR2_501(WX5036,WX5034,WX5033);
  or OR2_502(WX5043,WX5041,WX5040);
  or OR2_503(WX5050,WX5048,WX5047);
  or OR2_504(WX5057,WX5055,WX5054);
  or OR2_505(WX5064,WX5062,WX5061);
  or OR2_506(WX5071,WX5069,WX5068);
  or OR2_507(WX5078,WX5076,WX5075);
  or OR2_508(WX5085,WX5083,WX5082);
  or OR2_509(WX5092,WX5090,WX5089);
  or OR2_510(WX5099,WX5097,WX5096);
  or OR2_511(WX5106,WX5104,WX5103);
  or OR2_512(WX5210,WX5208,WX5207);
  or OR2_513(WX5214,WX5212,WX5211);
  or OR2_514(WX5218,WX5216,WX5215);
  or OR2_515(WX5224,WX5222,WX5221);
  or OR2_516(WX5228,WX5226,WX5225);
  or OR2_517(WX5232,WX5230,WX5229);
  or OR2_518(WX5238,WX5236,WX5235);
  or OR2_519(WX5242,WX5240,WX5239);
  or OR2_520(WX5246,WX5244,WX5243);
  or OR2_521(WX5252,WX5250,WX5249);
  or OR2_522(WX5256,WX5254,WX5253);
  or OR2_523(WX5260,WX5258,WX5257);
  or OR2_524(WX5266,WX5264,WX5263);
  or OR2_525(WX5270,WX5268,WX5267);
  or OR2_526(WX5274,WX5272,WX5271);
  or OR2_527(WX5280,WX5278,WX5277);
  or OR2_528(WX5284,WX5282,WX5281);
  or OR2_529(WX5288,WX5286,WX5285);
  or OR2_530(WX5294,WX5292,WX5291);
  or OR2_531(WX5298,WX5296,WX5295);
  or OR2_532(WX5302,WX5300,WX5299);
  or OR2_533(WX5308,WX5306,WX5305);
  or OR2_534(WX5312,WX5310,WX5309);
  or OR2_535(WX5316,WX5314,WX5313);
  or OR2_536(WX5322,WX5320,WX5319);
  or OR2_537(WX5326,WX5324,WX5323);
  or OR2_538(WX5330,WX5328,WX5327);
  or OR2_539(WX5336,WX5334,WX5333);
  or OR2_540(WX5340,WX5338,WX5337);
  or OR2_541(WX5344,WX5342,WX5341);
  or OR2_542(WX5350,WX5348,WX5347);
  or OR2_543(WX5354,WX5352,WX5351);
  or OR2_544(WX5358,WX5356,WX5355);
  or OR2_545(WX5364,WX5362,WX5361);
  or OR2_546(WX5368,WX5366,WX5365);
  or OR2_547(WX5372,WX5370,WX5369);
  or OR2_548(WX5378,WX5376,WX5375);
  or OR2_549(WX5382,WX5380,WX5379);
  or OR2_550(WX5386,WX5384,WX5383);
  or OR2_551(WX5392,WX5390,WX5389);
  or OR2_552(WX5396,WX5394,WX5393);
  or OR2_553(WX5400,WX5398,WX5397);
  or OR2_554(WX5406,WX5404,WX5403);
  or OR2_555(WX5410,WX5408,WX5407);
  or OR2_556(WX5414,WX5412,WX5411);
  or OR2_557(WX5420,WX5418,WX5417);
  or OR2_558(WX5424,WX5422,WX5421);
  or OR2_559(WX5428,WX5426,WX5425);
  or OR2_560(WX5434,WX5432,WX5431);
  or OR2_561(WX5438,WX5436,WX5435);
  or OR2_562(WX5442,WX5440,WX5439);
  or OR2_563(WX5448,WX5446,WX5445);
  or OR2_564(WX5452,WX5450,WX5449);
  or OR2_565(WX5456,WX5454,WX5453);
  or OR2_566(WX5462,WX5460,WX5459);
  or OR2_567(WX5466,WX5464,WX5463);
  or OR2_568(WX5470,WX5468,WX5467);
  or OR2_569(WX5476,WX5474,WX5473);
  or OR2_570(WX5480,WX5478,WX5477);
  or OR2_571(WX5484,WX5482,WX5481);
  or OR2_572(WX5490,WX5488,WX5487);
  or OR2_573(WX5494,WX5492,WX5491);
  or OR2_574(WX5498,WX5496,WX5495);
  or OR2_575(WX5504,WX5502,WX5501);
  or OR2_576(WX5508,WX5506,WX5505);
  or OR2_577(WX5512,WX5510,WX5509);
  or OR2_578(WX5518,WX5516,WX5515);
  or OR2_579(WX5522,WX5520,WX5519);
  or OR2_580(WX5526,WX5524,WX5523);
  or OR2_581(WX5532,WX5530,WX5529);
  or OR2_582(WX5536,WX5534,WX5533);
  or OR2_583(WX5540,WX5538,WX5537);
  or OR2_584(WX5546,WX5544,WX5543);
  or OR2_585(WX5550,WX5548,WX5547);
  or OR2_586(WX5554,WX5552,WX5551);
  or OR2_587(WX5560,WX5558,WX5557);
  or OR2_588(WX5564,WX5562,WX5561);
  or OR2_589(WX5568,WX5566,WX5565);
  or OR2_590(WX5574,WX5572,WX5571);
  or OR2_591(WX5578,WX5576,WX5575);
  or OR2_592(WX5582,WX5580,WX5579);
  or OR2_593(WX5588,WX5586,WX5585);
  or OR2_594(WX5592,WX5590,WX5589);
  or OR2_595(WX5596,WX5594,WX5593);
  or OR2_596(WX5602,WX5600,WX5599);
  or OR2_597(WX5606,WX5604,WX5603);
  or OR2_598(WX5610,WX5608,WX5607);
  or OR2_599(WX5616,WX5614,WX5613);
  or OR2_600(WX5620,WX5618,WX5617);
  or OR2_601(WX5624,WX5622,WX5621);
  or OR2_602(WX5630,WX5628,WX5627);
  or OR2_603(WX5634,WX5632,WX5631);
  or OR2_604(WX5638,WX5636,WX5635);
  or OR2_605(WX5644,WX5642,WX5641);
  or OR2_606(WX5648,WX5646,WX5645);
  or OR2_607(WX5652,WX5650,WX5649);
  or OR2_608(WX6182,WX6180,WX6179);
  or OR2_609(WX6189,WX6187,WX6186);
  or OR2_610(WX6196,WX6194,WX6193);
  or OR2_611(WX6203,WX6201,WX6200);
  or OR2_612(WX6210,WX6208,WX6207);
  or OR2_613(WX6217,WX6215,WX6214);
  or OR2_614(WX6224,WX6222,WX6221);
  or OR2_615(WX6231,WX6229,WX6228);
  or OR2_616(WX6238,WX6236,WX6235);
  or OR2_617(WX6245,WX6243,WX6242);
  or OR2_618(WX6252,WX6250,WX6249);
  or OR2_619(WX6259,WX6257,WX6256);
  or OR2_620(WX6266,WX6264,WX6263);
  or OR2_621(WX6273,WX6271,WX6270);
  or OR2_622(WX6280,WX6278,WX6277);
  or OR2_623(WX6287,WX6285,WX6284);
  or OR2_624(WX6294,WX6292,WX6291);
  or OR2_625(WX6301,WX6299,WX6298);
  or OR2_626(WX6308,WX6306,WX6305);
  or OR2_627(WX6315,WX6313,WX6312);
  or OR2_628(WX6322,WX6320,WX6319);
  or OR2_629(WX6329,WX6327,WX6326);
  or OR2_630(WX6336,WX6334,WX6333);
  or OR2_631(WX6343,WX6341,WX6340);
  or OR2_632(WX6350,WX6348,WX6347);
  or OR2_633(WX6357,WX6355,WX6354);
  or OR2_634(WX6364,WX6362,WX6361);
  or OR2_635(WX6371,WX6369,WX6368);
  or OR2_636(WX6378,WX6376,WX6375);
  or OR2_637(WX6385,WX6383,WX6382);
  or OR2_638(WX6392,WX6390,WX6389);
  or OR2_639(WX6399,WX6397,WX6396);
  or OR2_640(WX6503,WX6501,WX6500);
  or OR2_641(WX6507,WX6505,WX6504);
  or OR2_642(WX6511,WX6509,WX6508);
  or OR2_643(WX6517,WX6515,WX6514);
  or OR2_644(WX6521,WX6519,WX6518);
  or OR2_645(WX6525,WX6523,WX6522);
  or OR2_646(WX6531,WX6529,WX6528);
  or OR2_647(WX6535,WX6533,WX6532);
  or OR2_648(WX6539,WX6537,WX6536);
  or OR2_649(WX6545,WX6543,WX6542);
  or OR2_650(WX6549,WX6547,WX6546);
  or OR2_651(WX6553,WX6551,WX6550);
  or OR2_652(WX6559,WX6557,WX6556);
  or OR2_653(WX6563,WX6561,WX6560);
  or OR2_654(WX6567,WX6565,WX6564);
  or OR2_655(WX6573,WX6571,WX6570);
  or OR2_656(WX6577,WX6575,WX6574);
  or OR2_657(WX6581,WX6579,WX6578);
  or OR2_658(WX6587,WX6585,WX6584);
  or OR2_659(WX6591,WX6589,WX6588);
  or OR2_660(WX6595,WX6593,WX6592);
  or OR2_661(WX6601,WX6599,WX6598);
  or OR2_662(WX6605,WX6603,WX6602);
  or OR2_663(WX6609,WX6607,WX6606);
  or OR2_664(WX6615,WX6613,WX6612);
  or OR2_665(WX6619,WX6617,WX6616);
  or OR2_666(WX6623,WX6621,WX6620);
  or OR2_667(WX6629,WX6627,WX6626);
  or OR2_668(WX6633,WX6631,WX6630);
  or OR2_669(WX6637,WX6635,WX6634);
  or OR2_670(WX6643,WX6641,WX6640);
  or OR2_671(WX6647,WX6645,WX6644);
  or OR2_672(WX6651,WX6649,WX6648);
  or OR2_673(WX6657,WX6655,WX6654);
  or OR2_674(WX6661,WX6659,WX6658);
  or OR2_675(WX6665,WX6663,WX6662);
  or OR2_676(WX6671,WX6669,WX6668);
  or OR2_677(WX6675,WX6673,WX6672);
  or OR2_678(WX6679,WX6677,WX6676);
  or OR2_679(WX6685,WX6683,WX6682);
  or OR2_680(WX6689,WX6687,WX6686);
  or OR2_681(WX6693,WX6691,WX6690);
  or OR2_682(WX6699,WX6697,WX6696);
  or OR2_683(WX6703,WX6701,WX6700);
  or OR2_684(WX6707,WX6705,WX6704);
  or OR2_685(WX6713,WX6711,WX6710);
  or OR2_686(WX6717,WX6715,WX6714);
  or OR2_687(WX6721,WX6719,WX6718);
  or OR2_688(WX6727,WX6725,WX6724);
  or OR2_689(WX6731,WX6729,WX6728);
  or OR2_690(WX6735,WX6733,WX6732);
  or OR2_691(WX6741,WX6739,WX6738);
  or OR2_692(WX6745,WX6743,WX6742);
  or OR2_693(WX6749,WX6747,WX6746);
  or OR2_694(WX6755,WX6753,WX6752);
  or OR2_695(WX6759,WX6757,WX6756);
  or OR2_696(WX6763,WX6761,WX6760);
  or OR2_697(WX6769,WX6767,WX6766);
  or OR2_698(WX6773,WX6771,WX6770);
  or OR2_699(WX6777,WX6775,WX6774);
  or OR2_700(WX6783,WX6781,WX6780);
  or OR2_701(WX6787,WX6785,WX6784);
  or OR2_702(WX6791,WX6789,WX6788);
  or OR2_703(WX6797,WX6795,WX6794);
  or OR2_704(WX6801,WX6799,WX6798);
  or OR2_705(WX6805,WX6803,WX6802);
  or OR2_706(WX6811,WX6809,WX6808);
  or OR2_707(WX6815,WX6813,WX6812);
  or OR2_708(WX6819,WX6817,WX6816);
  or OR2_709(WX6825,WX6823,WX6822);
  or OR2_710(WX6829,WX6827,WX6826);
  or OR2_711(WX6833,WX6831,WX6830);
  or OR2_712(WX6839,WX6837,WX6836);
  or OR2_713(WX6843,WX6841,WX6840);
  or OR2_714(WX6847,WX6845,WX6844);
  or OR2_715(WX6853,WX6851,WX6850);
  or OR2_716(WX6857,WX6855,WX6854);
  or OR2_717(WX6861,WX6859,WX6858);
  or OR2_718(WX6867,WX6865,WX6864);
  or OR2_719(WX6871,WX6869,WX6868);
  or OR2_720(WX6875,WX6873,WX6872);
  or OR2_721(WX6881,WX6879,WX6878);
  or OR2_722(WX6885,WX6883,WX6882);
  or OR2_723(WX6889,WX6887,WX6886);
  or OR2_724(WX6895,WX6893,WX6892);
  or OR2_725(WX6899,WX6897,WX6896);
  or OR2_726(WX6903,WX6901,WX6900);
  or OR2_727(WX6909,WX6907,WX6906);
  or OR2_728(WX6913,WX6911,WX6910);
  or OR2_729(WX6917,WX6915,WX6914);
  or OR2_730(WX6923,WX6921,WX6920);
  or OR2_731(WX6927,WX6925,WX6924);
  or OR2_732(WX6931,WX6929,WX6928);
  or OR2_733(WX6937,WX6935,WX6934);
  or OR2_734(WX6941,WX6939,WX6938);
  or OR2_735(WX6945,WX6943,WX6942);
  or OR2_736(WX7475,WX7473,WX7472);
  or OR2_737(WX7482,WX7480,WX7479);
  or OR2_738(WX7489,WX7487,WX7486);
  or OR2_739(WX7496,WX7494,WX7493);
  or OR2_740(WX7503,WX7501,WX7500);
  or OR2_741(WX7510,WX7508,WX7507);
  or OR2_742(WX7517,WX7515,WX7514);
  or OR2_743(WX7524,WX7522,WX7521);
  or OR2_744(WX7531,WX7529,WX7528);
  or OR2_745(WX7538,WX7536,WX7535);
  or OR2_746(WX7545,WX7543,WX7542);
  or OR2_747(WX7552,WX7550,WX7549);
  or OR2_748(WX7559,WX7557,WX7556);
  or OR2_749(WX7566,WX7564,WX7563);
  or OR2_750(WX7573,WX7571,WX7570);
  or OR2_751(WX7580,WX7578,WX7577);
  or OR2_752(WX7587,WX7585,WX7584);
  or OR2_753(WX7594,WX7592,WX7591);
  or OR2_754(WX7601,WX7599,WX7598);
  or OR2_755(WX7608,WX7606,WX7605);
  or OR2_756(WX7615,WX7613,WX7612);
  or OR2_757(WX7622,WX7620,WX7619);
  or OR2_758(WX7629,WX7627,WX7626);
  or OR2_759(WX7636,WX7634,WX7633);
  or OR2_760(WX7643,WX7641,WX7640);
  or OR2_761(WX7650,WX7648,WX7647);
  or OR2_762(WX7657,WX7655,WX7654);
  or OR2_763(WX7664,WX7662,WX7661);
  or OR2_764(WX7671,WX7669,WX7668);
  or OR2_765(WX7678,WX7676,WX7675);
  or OR2_766(WX7685,WX7683,WX7682);
  or OR2_767(WX7692,WX7690,WX7689);
  or OR2_768(WX7796,WX7794,WX7793);
  or OR2_769(WX7800,WX7798,WX7797);
  or OR2_770(WX7804,WX7802,WX7801);
  or OR2_771(WX7810,WX7808,WX7807);
  or OR2_772(WX7814,WX7812,WX7811);
  or OR2_773(WX7818,WX7816,WX7815);
  or OR2_774(WX7824,WX7822,WX7821);
  or OR2_775(WX7828,WX7826,WX7825);
  or OR2_776(WX7832,WX7830,WX7829);
  or OR2_777(WX7838,WX7836,WX7835);
  or OR2_778(WX7842,WX7840,WX7839);
  or OR2_779(WX7846,WX7844,WX7843);
  or OR2_780(WX7852,WX7850,WX7849);
  or OR2_781(WX7856,WX7854,WX7853);
  or OR2_782(WX7860,WX7858,WX7857);
  or OR2_783(WX7866,WX7864,WX7863);
  or OR2_784(WX7870,WX7868,WX7867);
  or OR2_785(WX7874,WX7872,WX7871);
  or OR2_786(WX7880,WX7878,WX7877);
  or OR2_787(WX7884,WX7882,WX7881);
  or OR2_788(WX7888,WX7886,WX7885);
  or OR2_789(WX7894,WX7892,WX7891);
  or OR2_790(WX7898,WX7896,WX7895);
  or OR2_791(WX7902,WX7900,WX7899);
  or OR2_792(WX7908,WX7906,WX7905);
  or OR2_793(WX7912,WX7910,WX7909);
  or OR2_794(WX7916,WX7914,WX7913);
  or OR2_795(WX7922,WX7920,WX7919);
  or OR2_796(WX7926,WX7924,WX7923);
  or OR2_797(WX7930,WX7928,WX7927);
  or OR2_798(WX7936,WX7934,WX7933);
  or OR2_799(WX7940,WX7938,WX7937);
  or OR2_800(WX7944,WX7942,WX7941);
  or OR2_801(WX7950,WX7948,WX7947);
  or OR2_802(WX7954,WX7952,WX7951);
  or OR2_803(WX7958,WX7956,WX7955);
  or OR2_804(WX7964,WX7962,WX7961);
  or OR2_805(WX7968,WX7966,WX7965);
  or OR2_806(WX7972,WX7970,WX7969);
  or OR2_807(WX7978,WX7976,WX7975);
  or OR2_808(WX7982,WX7980,WX7979);
  or OR2_809(WX7986,WX7984,WX7983);
  or OR2_810(WX7992,WX7990,WX7989);
  or OR2_811(WX7996,WX7994,WX7993);
  or OR2_812(WX8000,WX7998,WX7997);
  or OR2_813(WX8006,WX8004,WX8003);
  or OR2_814(WX8010,WX8008,WX8007);
  or OR2_815(WX8014,WX8012,WX8011);
  or OR2_816(WX8020,WX8018,WX8017);
  or OR2_817(WX8024,WX8022,WX8021);
  or OR2_818(WX8028,WX8026,WX8025);
  or OR2_819(WX8034,WX8032,WX8031);
  or OR2_820(WX8038,WX8036,WX8035);
  or OR2_821(WX8042,WX8040,WX8039);
  or OR2_822(WX8048,WX8046,WX8045);
  or OR2_823(WX8052,WX8050,WX8049);
  or OR2_824(WX8056,WX8054,WX8053);
  or OR2_825(WX8062,WX8060,WX8059);
  or OR2_826(WX8066,WX8064,WX8063);
  or OR2_827(WX8070,WX8068,WX8067);
  or OR2_828(WX8076,WX8074,WX8073);
  or OR2_829(WX8080,WX8078,WX8077);
  or OR2_830(WX8084,WX8082,WX8081);
  or OR2_831(WX8090,WX8088,WX8087);
  or OR2_832(WX8094,WX8092,WX8091);
  or OR2_833(WX8098,WX8096,WX8095);
  or OR2_834(WX8104,WX8102,WX8101);
  or OR2_835(WX8108,WX8106,WX8105);
  or OR2_836(WX8112,WX8110,WX8109);
  or OR2_837(WX8118,WX8116,WX8115);
  or OR2_838(WX8122,WX8120,WX8119);
  or OR2_839(WX8126,WX8124,WX8123);
  or OR2_840(WX8132,WX8130,WX8129);
  or OR2_841(WX8136,WX8134,WX8133);
  or OR2_842(WX8140,WX8138,WX8137);
  or OR2_843(WX8146,WX8144,WX8143);
  or OR2_844(WX8150,WX8148,WX8147);
  or OR2_845(WX8154,WX8152,WX8151);
  or OR2_846(WX8160,WX8158,WX8157);
  or OR2_847(WX8164,WX8162,WX8161);
  or OR2_848(WX8168,WX8166,WX8165);
  or OR2_849(WX8174,WX8172,WX8171);
  or OR2_850(WX8178,WX8176,WX8175);
  or OR2_851(WX8182,WX8180,WX8179);
  or OR2_852(WX8188,WX8186,WX8185);
  or OR2_853(WX8192,WX8190,WX8189);
  or OR2_854(WX8196,WX8194,WX8193);
  or OR2_855(WX8202,WX8200,WX8199);
  or OR2_856(WX8206,WX8204,WX8203);
  or OR2_857(WX8210,WX8208,WX8207);
  or OR2_858(WX8216,WX8214,WX8213);
  or OR2_859(WX8220,WX8218,WX8217);
  or OR2_860(WX8224,WX8222,WX8221);
  or OR2_861(WX8230,WX8228,WX8227);
  or OR2_862(WX8234,WX8232,WX8231);
  or OR2_863(WX8238,WX8236,WX8235);
  or OR2_864(WX8768,WX8766,WX8765);
  or OR2_865(WX8775,WX8773,WX8772);
  or OR2_866(WX8782,WX8780,WX8779);
  or OR2_867(WX8789,WX8787,WX8786);
  or OR2_868(WX8796,WX8794,WX8793);
  or OR2_869(WX8803,WX8801,WX8800);
  or OR2_870(WX8810,WX8808,WX8807);
  or OR2_871(WX8817,WX8815,WX8814);
  or OR2_872(WX8824,WX8822,WX8821);
  or OR2_873(WX8831,WX8829,WX8828);
  or OR2_874(WX8838,WX8836,WX8835);
  or OR2_875(WX8845,WX8843,WX8842);
  or OR2_876(WX8852,WX8850,WX8849);
  or OR2_877(WX8859,WX8857,WX8856);
  or OR2_878(WX8866,WX8864,WX8863);
  or OR2_879(WX8873,WX8871,WX8870);
  or OR2_880(WX8880,WX8878,WX8877);
  or OR2_881(WX8887,WX8885,WX8884);
  or OR2_882(WX8894,WX8892,WX8891);
  or OR2_883(WX8901,WX8899,WX8898);
  or OR2_884(WX8908,WX8906,WX8905);
  or OR2_885(WX8915,WX8913,WX8912);
  or OR2_886(WX8922,WX8920,WX8919);
  or OR2_887(WX8929,WX8927,WX8926);
  or OR2_888(WX8936,WX8934,WX8933);
  or OR2_889(WX8943,WX8941,WX8940);
  or OR2_890(WX8950,WX8948,WX8947);
  or OR2_891(WX8957,WX8955,WX8954);
  or OR2_892(WX8964,WX8962,WX8961);
  or OR2_893(WX8971,WX8969,WX8968);
  or OR2_894(WX8978,WX8976,WX8975);
  or OR2_895(WX8985,WX8983,WX8982);
  or OR2_896(WX9089,WX9087,WX9086);
  or OR2_897(WX9093,WX9091,WX9090);
  or OR2_898(WX9097,WX9095,WX9094);
  or OR2_899(WX9103,WX9101,WX9100);
  or OR2_900(WX9107,WX9105,WX9104);
  or OR2_901(WX9111,WX9109,WX9108);
  or OR2_902(WX9117,WX9115,WX9114);
  or OR2_903(WX9121,WX9119,WX9118);
  or OR2_904(WX9125,WX9123,WX9122);
  or OR2_905(WX9131,WX9129,WX9128);
  or OR2_906(WX9135,WX9133,WX9132);
  or OR2_907(WX9139,WX9137,WX9136);
  or OR2_908(WX9145,WX9143,WX9142);
  or OR2_909(WX9149,WX9147,WX9146);
  or OR2_910(WX9153,WX9151,WX9150);
  or OR2_911(WX9159,WX9157,WX9156);
  or OR2_912(WX9163,WX9161,WX9160);
  or OR2_913(WX9167,WX9165,WX9164);
  or OR2_914(WX9173,WX9171,WX9170);
  or OR2_915(WX9177,WX9175,WX9174);
  or OR2_916(WX9181,WX9179,WX9178);
  or OR2_917(WX9187,WX9185,WX9184);
  or OR2_918(WX9191,WX9189,WX9188);
  or OR2_919(WX9195,WX9193,WX9192);
  or OR2_920(WX9201,WX9199,WX9198);
  or OR2_921(WX9205,WX9203,WX9202);
  or OR2_922(WX9209,WX9207,WX9206);
  or OR2_923(WX9215,WX9213,WX9212);
  or OR2_924(WX9219,WX9217,WX9216);
  or OR2_925(WX9223,WX9221,WX9220);
  or OR2_926(WX9229,WX9227,WX9226);
  or OR2_927(WX9233,WX9231,WX9230);
  or OR2_928(WX9237,WX9235,WX9234);
  or OR2_929(WX9243,WX9241,WX9240);
  or OR2_930(WX9247,WX9245,WX9244);
  or OR2_931(WX9251,WX9249,WX9248);
  or OR2_932(WX9257,WX9255,WX9254);
  or OR2_933(WX9261,WX9259,WX9258);
  or OR2_934(WX9265,WX9263,WX9262);
  or OR2_935(WX9271,WX9269,WX9268);
  or OR2_936(WX9275,WX9273,WX9272);
  or OR2_937(WX9279,WX9277,WX9276);
  or OR2_938(WX9285,WX9283,WX9282);
  or OR2_939(WX9289,WX9287,WX9286);
  or OR2_940(WX9293,WX9291,WX9290);
  or OR2_941(WX9299,WX9297,WX9296);
  or OR2_942(WX9303,WX9301,WX9300);
  or OR2_943(WX9307,WX9305,WX9304);
  or OR2_944(WX9313,WX9311,WX9310);
  or OR2_945(WX9317,WX9315,WX9314);
  or OR2_946(WX9321,WX9319,WX9318);
  or OR2_947(WX9327,WX9325,WX9324);
  or OR2_948(WX9331,WX9329,WX9328);
  or OR2_949(WX9335,WX9333,WX9332);
  or OR2_950(WX9341,WX9339,WX9338);
  or OR2_951(WX9345,WX9343,WX9342);
  or OR2_952(WX9349,WX9347,WX9346);
  or OR2_953(WX9355,WX9353,WX9352);
  or OR2_954(WX9359,WX9357,WX9356);
  or OR2_955(WX9363,WX9361,WX9360);
  or OR2_956(WX9369,WX9367,WX9366);
  or OR2_957(WX9373,WX9371,WX9370);
  or OR2_958(WX9377,WX9375,WX9374);
  or OR2_959(WX9383,WX9381,WX9380);
  or OR2_960(WX9387,WX9385,WX9384);
  or OR2_961(WX9391,WX9389,WX9388);
  or OR2_962(WX9397,WX9395,WX9394);
  or OR2_963(WX9401,WX9399,WX9398);
  or OR2_964(WX9405,WX9403,WX9402);
  or OR2_965(WX9411,WX9409,WX9408);
  or OR2_966(WX9415,WX9413,WX9412);
  or OR2_967(WX9419,WX9417,WX9416);
  or OR2_968(WX9425,WX9423,WX9422);
  or OR2_969(WX9429,WX9427,WX9426);
  or OR2_970(WX9433,WX9431,WX9430);
  or OR2_971(WX9439,WX9437,WX9436);
  or OR2_972(WX9443,WX9441,WX9440);
  or OR2_973(WX9447,WX9445,WX9444);
  or OR2_974(WX9453,WX9451,WX9450);
  or OR2_975(WX9457,WX9455,WX9454);
  or OR2_976(WX9461,WX9459,WX9458);
  or OR2_977(WX9467,WX9465,WX9464);
  or OR2_978(WX9471,WX9469,WX9468);
  or OR2_979(WX9475,WX9473,WX9472);
  or OR2_980(WX9481,WX9479,WX9478);
  or OR2_981(WX9485,WX9483,WX9482);
  or OR2_982(WX9489,WX9487,WX9486);
  or OR2_983(WX9495,WX9493,WX9492);
  or OR2_984(WX9499,WX9497,WX9496);
  or OR2_985(WX9503,WX9501,WX9500);
  or OR2_986(WX9509,WX9507,WX9506);
  or OR2_987(WX9513,WX9511,WX9510);
  or OR2_988(WX9517,WX9515,WX9514);
  or OR2_989(WX9523,WX9521,WX9520);
  or OR2_990(WX9527,WX9525,WX9524);
  or OR2_991(WX9531,WX9529,WX9528);
  or OR2_992(WX10061,WX10059,WX10058);
  or OR2_993(WX10068,WX10066,WX10065);
  or OR2_994(WX10075,WX10073,WX10072);
  or OR2_995(WX10082,WX10080,WX10079);
  or OR2_996(WX10089,WX10087,WX10086);
  or OR2_997(WX10096,WX10094,WX10093);
  or OR2_998(WX10103,WX10101,WX10100);
  or OR2_999(WX10110,WX10108,WX10107);
  or OR2_1000(WX10117,WX10115,WX10114);
  or OR2_1001(WX10124,WX10122,WX10121);
  or OR2_1002(WX10131,WX10129,WX10128);
  or OR2_1003(WX10138,WX10136,WX10135);
  or OR2_1004(WX10145,WX10143,WX10142);
  or OR2_1005(WX10152,WX10150,WX10149);
  or OR2_1006(WX10159,WX10157,WX10156);
  or OR2_1007(WX10166,WX10164,WX10163);
  or OR2_1008(WX10173,WX10171,WX10170);
  or OR2_1009(WX10180,WX10178,WX10177);
  or OR2_1010(WX10187,WX10185,WX10184);
  or OR2_1011(WX10194,WX10192,WX10191);
  or OR2_1012(WX10201,WX10199,WX10198);
  or OR2_1013(WX10208,WX10206,WX10205);
  or OR2_1014(WX10215,WX10213,WX10212);
  or OR2_1015(WX10222,WX10220,WX10219);
  or OR2_1016(WX10229,WX10227,WX10226);
  or OR2_1017(WX10236,WX10234,WX10233);
  or OR2_1018(WX10243,WX10241,WX10240);
  or OR2_1019(WX10250,WX10248,WX10247);
  or OR2_1020(WX10257,WX10255,WX10254);
  or OR2_1021(WX10264,WX10262,WX10261);
  or OR2_1022(WX10271,WX10269,WX10268);
  or OR2_1023(WX10278,WX10276,WX10275);
  or OR2_1024(WX10382,WX10380,WX10379);
  or OR2_1025(WX10386,WX10384,WX10383);
  or OR2_1026(WX10390,WX10388,WX10387);
  or OR2_1027(WX10396,WX10394,WX10393);
  or OR2_1028(WX10400,WX10398,WX10397);
  or OR2_1029(WX10404,WX10402,WX10401);
  or OR2_1030(WX10410,WX10408,WX10407);
  or OR2_1031(WX10414,WX10412,WX10411);
  or OR2_1032(WX10418,WX10416,WX10415);
  or OR2_1033(WX10424,WX10422,WX10421);
  or OR2_1034(WX10428,WX10426,WX10425);
  or OR2_1035(WX10432,WX10430,WX10429);
  or OR2_1036(WX10438,WX10436,WX10435);
  or OR2_1037(WX10442,WX10440,WX10439);
  or OR2_1038(WX10446,WX10444,WX10443);
  or OR2_1039(WX10452,WX10450,WX10449);
  or OR2_1040(WX10456,WX10454,WX10453);
  or OR2_1041(WX10460,WX10458,WX10457);
  or OR2_1042(WX10466,WX10464,WX10463);
  or OR2_1043(WX10470,WX10468,WX10467);
  or OR2_1044(WX10474,WX10472,WX10471);
  or OR2_1045(WX10480,WX10478,WX10477);
  or OR2_1046(WX10484,WX10482,WX10481);
  or OR2_1047(WX10488,WX10486,WX10485);
  or OR2_1048(WX10494,WX10492,WX10491);
  or OR2_1049(WX10498,WX10496,WX10495);
  or OR2_1050(WX10502,WX10500,WX10499);
  or OR2_1051(WX10508,WX10506,WX10505);
  or OR2_1052(WX10512,WX10510,WX10509);
  or OR2_1053(WX10516,WX10514,WX10513);
  or OR2_1054(WX10522,WX10520,WX10519);
  or OR2_1055(WX10526,WX10524,WX10523);
  or OR2_1056(WX10530,WX10528,WX10527);
  or OR2_1057(WX10536,WX10534,WX10533);
  or OR2_1058(WX10540,WX10538,WX10537);
  or OR2_1059(WX10544,WX10542,WX10541);
  or OR2_1060(WX10550,WX10548,WX10547);
  or OR2_1061(WX10554,WX10552,WX10551);
  or OR2_1062(WX10558,WX10556,WX10555);
  or OR2_1063(WX10564,WX10562,WX10561);
  or OR2_1064(WX10568,WX10566,WX10565);
  or OR2_1065(WX10572,WX10570,WX10569);
  or OR2_1066(WX10578,WX10576,WX10575);
  or OR2_1067(WX10582,WX10580,WX10579);
  or OR2_1068(WX10586,WX10584,WX10583);
  or OR2_1069(WX10592,WX10590,WX10589);
  or OR2_1070(WX10596,WX10594,WX10593);
  or OR2_1071(WX10600,WX10598,WX10597);
  or OR2_1072(WX10606,WX10604,WX10603);
  or OR2_1073(WX10610,WX10608,WX10607);
  or OR2_1074(WX10614,WX10612,WX10611);
  or OR2_1075(WX10620,WX10618,WX10617);
  or OR2_1076(WX10624,WX10622,WX10621);
  or OR2_1077(WX10628,WX10626,WX10625);
  or OR2_1078(WX10634,WX10632,WX10631);
  or OR2_1079(WX10638,WX10636,WX10635);
  or OR2_1080(WX10642,WX10640,WX10639);
  or OR2_1081(WX10648,WX10646,WX10645);
  or OR2_1082(WX10652,WX10650,WX10649);
  or OR2_1083(WX10656,WX10654,WX10653);
  or OR2_1084(WX10662,WX10660,WX10659);
  or OR2_1085(WX10666,WX10664,WX10663);
  or OR2_1086(WX10670,WX10668,WX10667);
  or OR2_1087(WX10676,WX10674,WX10673);
  or OR2_1088(WX10680,WX10678,WX10677);
  or OR2_1089(WX10684,WX10682,WX10681);
  or OR2_1090(WX10690,WX10688,WX10687);
  or OR2_1091(WX10694,WX10692,WX10691);
  or OR2_1092(WX10698,WX10696,WX10695);
  or OR2_1093(WX10704,WX10702,WX10701);
  or OR2_1094(WX10708,WX10706,WX10705);
  or OR2_1095(WX10712,WX10710,WX10709);
  or OR2_1096(WX10718,WX10716,WX10715);
  or OR2_1097(WX10722,WX10720,WX10719);
  or OR2_1098(WX10726,WX10724,WX10723);
  or OR2_1099(WX10732,WX10730,WX10729);
  or OR2_1100(WX10736,WX10734,WX10733);
  or OR2_1101(WX10740,WX10738,WX10737);
  or OR2_1102(WX10746,WX10744,WX10743);
  or OR2_1103(WX10750,WX10748,WX10747);
  or OR2_1104(WX10754,WX10752,WX10751);
  or OR2_1105(WX10760,WX10758,WX10757);
  or OR2_1106(WX10764,WX10762,WX10761);
  or OR2_1107(WX10768,WX10766,WX10765);
  or OR2_1108(WX10774,WX10772,WX10771);
  or OR2_1109(WX10778,WX10776,WX10775);
  or OR2_1110(WX10782,WX10780,WX10779);
  or OR2_1111(WX10788,WX10786,WX10785);
  or OR2_1112(WX10792,WX10790,WX10789);
  or OR2_1113(WX10796,WX10794,WX10793);
  or OR2_1114(WX10802,WX10800,WX10799);
  or OR2_1115(WX10806,WX10804,WX10803);
  or OR2_1116(WX10810,WX10808,WX10807);
  or OR2_1117(WX10816,WX10814,WX10813);
  or OR2_1118(WX10820,WX10818,WX10817);
  or OR2_1119(WX10824,WX10822,WX10821);
  or OR2_1120(WX11354,WX11352,WX11351);
  or OR2_1121(WX11361,WX11359,WX11358);
  or OR2_1122(WX11368,WX11366,WX11365);
  or OR2_1123(WX11375,WX11373,WX11372);
  or OR2_1124(WX11382,WX11380,WX11379);
  or OR2_1125(WX11389,WX11387,WX11386);
  or OR2_1126(WX11396,WX11394,WX11393);
  or OR2_1127(WX11403,WX11401,WX11400);
  or OR2_1128(WX11410,WX11408,WX11407);
  or OR2_1129(WX11417,WX11415,WX11414);
  or OR2_1130(WX11424,WX11422,WX11421);
  or OR2_1131(WX11431,WX11429,WX11428);
  or OR2_1132(WX11438,WX11436,WX11435);
  or OR2_1133(WX11445,WX11443,WX11442);
  or OR2_1134(WX11452,WX11450,WX11449);
  or OR2_1135(WX11459,WX11457,WX11456);
  or OR2_1136(WX11466,WX11464,WX11463);
  or OR2_1137(WX11473,WX11471,WX11470);
  or OR2_1138(WX11480,WX11478,WX11477);
  or OR2_1139(WX11487,WX11485,WX11484);
  or OR2_1140(WX11494,WX11492,WX11491);
  or OR2_1141(WX11501,WX11499,WX11498);
  or OR2_1142(WX11508,WX11506,WX11505);
  or OR2_1143(WX11515,WX11513,WX11512);
  or OR2_1144(WX11522,WX11520,WX11519);
  or OR2_1145(WX11529,WX11527,WX11526);
  or OR2_1146(WX11536,WX11534,WX11533);
  or OR2_1147(WX11543,WX11541,WX11540);
  or OR2_1148(WX11550,WX11548,WX11547);
  or OR2_1149(WX11557,WX11555,WX11554);
  or OR2_1150(WX11564,WX11562,WX11561);
  or OR2_1151(WX11571,WX11569,WX11568);
  nand NAND2_0(II1988,WX1001,WX645);
  nand NAND2_1(II1989,WX1001,II1988);
  nand NAND2_2(II1990,WX645,II1988);
  nand NAND2_3(II1987,II1989,II1990);
  nand NAND2_4(II1995,WX709,II1987);
  nand NAND2_5(II1996,WX709,II1995);
  nand NAND2_6(II1997,II1987,II1995);
  nand NAND2_7(II1986,II1996,II1997);
  nand NAND2_8(II2003,WX773,WX837);
  nand NAND2_9(II2004,WX773,II2003);
  nand NAND2_10(II2005,WX837,II2003);
  nand NAND2_11(II2002,II2004,II2005);
  nand NAND2_12(II2010,II1986,II2002);
  nand NAND2_13(II2011,II1986,II2010);
  nand NAND2_14(II2012,II2002,II2010);
  nand NAND2_15(WX900,II2011,II2012);
  nand NAND2_16(II2019,WX1001,WX647);
  nand NAND2_17(II2020,WX1001,II2019);
  nand NAND2_18(II2021,WX647,II2019);
  nand NAND2_19(II2018,II2020,II2021);
  nand NAND2_20(II2026,WX711,II2018);
  nand NAND2_21(II2027,WX711,II2026);
  nand NAND2_22(II2028,II2018,II2026);
  nand NAND2_23(II2017,II2027,II2028);
  nand NAND2_24(II2034,WX775,WX839);
  nand NAND2_25(II2035,WX775,II2034);
  nand NAND2_26(II2036,WX839,II2034);
  nand NAND2_27(II2033,II2035,II2036);
  nand NAND2_28(II2041,II2017,II2033);
  nand NAND2_29(II2042,II2017,II2041);
  nand NAND2_30(II2043,II2033,II2041);
  nand NAND2_31(WX901,II2042,II2043);
  nand NAND2_32(II2050,WX1001,WX649);
  nand NAND2_33(II2051,WX1001,II2050);
  nand NAND2_34(II2052,WX649,II2050);
  nand NAND2_35(II2049,II2051,II2052);
  nand NAND2_36(II2057,WX713,II2049);
  nand NAND2_37(II2058,WX713,II2057);
  nand NAND2_38(II2059,II2049,II2057);
  nand NAND2_39(II2048,II2058,II2059);
  nand NAND2_40(II2065,WX777,WX841);
  nand NAND2_41(II2066,WX777,II2065);
  nand NAND2_42(II2067,WX841,II2065);
  nand NAND2_43(II2064,II2066,II2067);
  nand NAND2_44(II2072,II2048,II2064);
  nand NAND2_45(II2073,II2048,II2072);
  nand NAND2_46(II2074,II2064,II2072);
  nand NAND2_47(WX902,II2073,II2074);
  nand NAND2_48(II2081,WX1001,WX651);
  nand NAND2_49(II2082,WX1001,II2081);
  nand NAND2_50(II2083,WX651,II2081);
  nand NAND2_51(II2080,II2082,II2083);
  nand NAND2_52(II2088,WX715,II2080);
  nand NAND2_53(II2089,WX715,II2088);
  nand NAND2_54(II2090,II2080,II2088);
  nand NAND2_55(II2079,II2089,II2090);
  nand NAND2_56(II2096,WX779,WX843);
  nand NAND2_57(II2097,WX779,II2096);
  nand NAND2_58(II2098,WX843,II2096);
  nand NAND2_59(II2095,II2097,II2098);
  nand NAND2_60(II2103,II2079,II2095);
  nand NAND2_61(II2104,II2079,II2103);
  nand NAND2_62(II2105,II2095,II2103);
  nand NAND2_63(WX903,II2104,II2105);
  nand NAND2_64(II2112,WX1001,WX653);
  nand NAND2_65(II2113,WX1001,II2112);
  nand NAND2_66(II2114,WX653,II2112);
  nand NAND2_67(II2111,II2113,II2114);
  nand NAND2_68(II2119,WX717,II2111);
  nand NAND2_69(II2120,WX717,II2119);
  nand NAND2_70(II2121,II2111,II2119);
  nand NAND2_71(II2110,II2120,II2121);
  nand NAND2_72(II2127,WX781,WX845);
  nand NAND2_73(II2128,WX781,II2127);
  nand NAND2_74(II2129,WX845,II2127);
  nand NAND2_75(II2126,II2128,II2129);
  nand NAND2_76(II2134,II2110,II2126);
  nand NAND2_77(II2135,II2110,II2134);
  nand NAND2_78(II2136,II2126,II2134);
  nand NAND2_79(WX904,II2135,II2136);
  nand NAND2_80(II2143,WX1001,WX655);
  nand NAND2_81(II2144,WX1001,II2143);
  nand NAND2_82(II2145,WX655,II2143);
  nand NAND2_83(II2142,II2144,II2145);
  nand NAND2_84(II2150,WX719,II2142);
  nand NAND2_85(II2151,WX719,II2150);
  nand NAND2_86(II2152,II2142,II2150);
  nand NAND2_87(II2141,II2151,II2152);
  nand NAND2_88(II2158,WX783,WX847);
  nand NAND2_89(II2159,WX783,II2158);
  nand NAND2_90(II2160,WX847,II2158);
  nand NAND2_91(II2157,II2159,II2160);
  nand NAND2_92(II2165,II2141,II2157);
  nand NAND2_93(II2166,II2141,II2165);
  nand NAND2_94(II2167,II2157,II2165);
  nand NAND2_95(WX905,II2166,II2167);
  nand NAND2_96(II2174,WX1001,WX657);
  nand NAND2_97(II2175,WX1001,II2174);
  nand NAND2_98(II2176,WX657,II2174);
  nand NAND2_99(II2173,II2175,II2176);
  nand NAND2_100(II2181,WX721,II2173);
  nand NAND2_101(II2182,WX721,II2181);
  nand NAND2_102(II2183,II2173,II2181);
  nand NAND2_103(II2172,II2182,II2183);
  nand NAND2_104(II2189,WX785,WX849);
  nand NAND2_105(II2190,WX785,II2189);
  nand NAND2_106(II2191,WX849,II2189);
  nand NAND2_107(II2188,II2190,II2191);
  nand NAND2_108(II2196,II2172,II2188);
  nand NAND2_109(II2197,II2172,II2196);
  nand NAND2_110(II2198,II2188,II2196);
  nand NAND2_111(WX906,II2197,II2198);
  nand NAND2_112(II2205,WX1001,WX659);
  nand NAND2_113(II2206,WX1001,II2205);
  nand NAND2_114(II2207,WX659,II2205);
  nand NAND2_115(II2204,II2206,II2207);
  nand NAND2_116(II2212,WX723,II2204);
  nand NAND2_117(II2213,WX723,II2212);
  nand NAND2_118(II2214,II2204,II2212);
  nand NAND2_119(II2203,II2213,II2214);
  nand NAND2_120(II2220,WX787,WX851);
  nand NAND2_121(II2221,WX787,II2220);
  nand NAND2_122(II2222,WX851,II2220);
  nand NAND2_123(II2219,II2221,II2222);
  nand NAND2_124(II2227,II2203,II2219);
  nand NAND2_125(II2228,II2203,II2227);
  nand NAND2_126(II2229,II2219,II2227);
  nand NAND2_127(WX907,II2228,II2229);
  nand NAND2_128(II2236,WX1001,WX661);
  nand NAND2_129(II2237,WX1001,II2236);
  nand NAND2_130(II2238,WX661,II2236);
  nand NAND2_131(II2235,II2237,II2238);
  nand NAND2_132(II2243,WX725,II2235);
  nand NAND2_133(II2244,WX725,II2243);
  nand NAND2_134(II2245,II2235,II2243);
  nand NAND2_135(II2234,II2244,II2245);
  nand NAND2_136(II2251,WX789,WX853);
  nand NAND2_137(II2252,WX789,II2251);
  nand NAND2_138(II2253,WX853,II2251);
  nand NAND2_139(II2250,II2252,II2253);
  nand NAND2_140(II2258,II2234,II2250);
  nand NAND2_141(II2259,II2234,II2258);
  nand NAND2_142(II2260,II2250,II2258);
  nand NAND2_143(WX908,II2259,II2260);
  nand NAND2_144(II2267,WX1001,WX663);
  nand NAND2_145(II2268,WX1001,II2267);
  nand NAND2_146(II2269,WX663,II2267);
  nand NAND2_147(II2266,II2268,II2269);
  nand NAND2_148(II2274,WX727,II2266);
  nand NAND2_149(II2275,WX727,II2274);
  nand NAND2_150(II2276,II2266,II2274);
  nand NAND2_151(II2265,II2275,II2276);
  nand NAND2_152(II2282,WX791,WX855);
  nand NAND2_153(II2283,WX791,II2282);
  nand NAND2_154(II2284,WX855,II2282);
  nand NAND2_155(II2281,II2283,II2284);
  nand NAND2_156(II2289,II2265,II2281);
  nand NAND2_157(II2290,II2265,II2289);
  nand NAND2_158(II2291,II2281,II2289);
  nand NAND2_159(WX909,II2290,II2291);
  nand NAND2_160(II2298,WX1001,WX665);
  nand NAND2_161(II2299,WX1001,II2298);
  nand NAND2_162(II2300,WX665,II2298);
  nand NAND2_163(II2297,II2299,II2300);
  nand NAND2_164(II2305,WX729,II2297);
  nand NAND2_165(II2306,WX729,II2305);
  nand NAND2_166(II2307,II2297,II2305);
  nand NAND2_167(II2296,II2306,II2307);
  nand NAND2_168(II2313,WX793,WX857);
  nand NAND2_169(II2314,WX793,II2313);
  nand NAND2_170(II2315,WX857,II2313);
  nand NAND2_171(II2312,II2314,II2315);
  nand NAND2_172(II2320,II2296,II2312);
  nand NAND2_173(II2321,II2296,II2320);
  nand NAND2_174(II2322,II2312,II2320);
  nand NAND2_175(WX910,II2321,II2322);
  nand NAND2_176(II2329,WX1001,WX667);
  nand NAND2_177(II2330,WX1001,II2329);
  nand NAND2_178(II2331,WX667,II2329);
  nand NAND2_179(II2328,II2330,II2331);
  nand NAND2_180(II2336,WX731,II2328);
  nand NAND2_181(II2337,WX731,II2336);
  nand NAND2_182(II2338,II2328,II2336);
  nand NAND2_183(II2327,II2337,II2338);
  nand NAND2_184(II2344,WX795,WX859);
  nand NAND2_185(II2345,WX795,II2344);
  nand NAND2_186(II2346,WX859,II2344);
  nand NAND2_187(II2343,II2345,II2346);
  nand NAND2_188(II2351,II2327,II2343);
  nand NAND2_189(II2352,II2327,II2351);
  nand NAND2_190(II2353,II2343,II2351);
  nand NAND2_191(WX911,II2352,II2353);
  nand NAND2_192(II2360,WX1001,WX669);
  nand NAND2_193(II2361,WX1001,II2360);
  nand NAND2_194(II2362,WX669,II2360);
  nand NAND2_195(II2359,II2361,II2362);
  nand NAND2_196(II2367,WX733,II2359);
  nand NAND2_197(II2368,WX733,II2367);
  nand NAND2_198(II2369,II2359,II2367);
  nand NAND2_199(II2358,II2368,II2369);
  nand NAND2_200(II2375,WX797,WX861);
  nand NAND2_201(II2376,WX797,II2375);
  nand NAND2_202(II2377,WX861,II2375);
  nand NAND2_203(II2374,II2376,II2377);
  nand NAND2_204(II2382,II2358,II2374);
  nand NAND2_205(II2383,II2358,II2382);
  nand NAND2_206(II2384,II2374,II2382);
  nand NAND2_207(WX912,II2383,II2384);
  nand NAND2_208(II2391,WX1001,WX671);
  nand NAND2_209(II2392,WX1001,II2391);
  nand NAND2_210(II2393,WX671,II2391);
  nand NAND2_211(II2390,II2392,II2393);
  nand NAND2_212(II2398,WX735,II2390);
  nand NAND2_213(II2399,WX735,II2398);
  nand NAND2_214(II2400,II2390,II2398);
  nand NAND2_215(II2389,II2399,II2400);
  nand NAND2_216(II2406,WX799,WX863);
  nand NAND2_217(II2407,WX799,II2406);
  nand NAND2_218(II2408,WX863,II2406);
  nand NAND2_219(II2405,II2407,II2408);
  nand NAND2_220(II2413,II2389,II2405);
  nand NAND2_221(II2414,II2389,II2413);
  nand NAND2_222(II2415,II2405,II2413);
  nand NAND2_223(WX913,II2414,II2415);
  nand NAND2_224(II2422,WX1001,WX673);
  nand NAND2_225(II2423,WX1001,II2422);
  nand NAND2_226(II2424,WX673,II2422);
  nand NAND2_227(II2421,II2423,II2424);
  nand NAND2_228(II2429,WX737,II2421);
  nand NAND2_229(II2430,WX737,II2429);
  nand NAND2_230(II2431,II2421,II2429);
  nand NAND2_231(II2420,II2430,II2431);
  nand NAND2_232(II2437,WX801,WX865);
  nand NAND2_233(II2438,WX801,II2437);
  nand NAND2_234(II2439,WX865,II2437);
  nand NAND2_235(II2436,II2438,II2439);
  nand NAND2_236(II2444,II2420,II2436);
  nand NAND2_237(II2445,II2420,II2444);
  nand NAND2_238(II2446,II2436,II2444);
  nand NAND2_239(WX914,II2445,II2446);
  nand NAND2_240(II2453,WX1001,WX675);
  nand NAND2_241(II2454,WX1001,II2453);
  nand NAND2_242(II2455,WX675,II2453);
  nand NAND2_243(II2452,II2454,II2455);
  nand NAND2_244(II2460,WX739,II2452);
  nand NAND2_245(II2461,WX739,II2460);
  nand NAND2_246(II2462,II2452,II2460);
  nand NAND2_247(II2451,II2461,II2462);
  nand NAND2_248(II2468,WX803,WX867);
  nand NAND2_249(II2469,WX803,II2468);
  nand NAND2_250(II2470,WX867,II2468);
  nand NAND2_251(II2467,II2469,II2470);
  nand NAND2_252(II2475,II2451,II2467);
  nand NAND2_253(II2476,II2451,II2475);
  nand NAND2_254(II2477,II2467,II2475);
  nand NAND2_255(WX915,II2476,II2477);
  nand NAND2_256(II2484,WX1002,WX677);
  nand NAND2_257(II2485,WX1002,II2484);
  nand NAND2_258(II2486,WX677,II2484);
  nand NAND2_259(II2483,II2485,II2486);
  nand NAND2_260(II2491,WX741,II2483);
  nand NAND2_261(II2492,WX741,II2491);
  nand NAND2_262(II2493,II2483,II2491);
  nand NAND2_263(II2482,II2492,II2493);
  nand NAND2_264(II2499,WX805,WX869);
  nand NAND2_265(II2500,WX805,II2499);
  nand NAND2_266(II2501,WX869,II2499);
  nand NAND2_267(II2498,II2500,II2501);
  nand NAND2_268(II2506,II2482,II2498);
  nand NAND2_269(II2507,II2482,II2506);
  nand NAND2_270(II2508,II2498,II2506);
  nand NAND2_271(WX916,II2507,II2508);
  nand NAND2_272(II2515,WX1002,WX679);
  nand NAND2_273(II2516,WX1002,II2515);
  nand NAND2_274(II2517,WX679,II2515);
  nand NAND2_275(II2514,II2516,II2517);
  nand NAND2_276(II2522,WX743,II2514);
  nand NAND2_277(II2523,WX743,II2522);
  nand NAND2_278(II2524,II2514,II2522);
  nand NAND2_279(II2513,II2523,II2524);
  nand NAND2_280(II2530,WX807,WX871);
  nand NAND2_281(II2531,WX807,II2530);
  nand NAND2_282(II2532,WX871,II2530);
  nand NAND2_283(II2529,II2531,II2532);
  nand NAND2_284(II2537,II2513,II2529);
  nand NAND2_285(II2538,II2513,II2537);
  nand NAND2_286(II2539,II2529,II2537);
  nand NAND2_287(WX917,II2538,II2539);
  nand NAND2_288(II2546,WX1002,WX681);
  nand NAND2_289(II2547,WX1002,II2546);
  nand NAND2_290(II2548,WX681,II2546);
  nand NAND2_291(II2545,II2547,II2548);
  nand NAND2_292(II2553,WX745,II2545);
  nand NAND2_293(II2554,WX745,II2553);
  nand NAND2_294(II2555,II2545,II2553);
  nand NAND2_295(II2544,II2554,II2555);
  nand NAND2_296(II2561,WX809,WX873);
  nand NAND2_297(II2562,WX809,II2561);
  nand NAND2_298(II2563,WX873,II2561);
  nand NAND2_299(II2560,II2562,II2563);
  nand NAND2_300(II2568,II2544,II2560);
  nand NAND2_301(II2569,II2544,II2568);
  nand NAND2_302(II2570,II2560,II2568);
  nand NAND2_303(WX918,II2569,II2570);
  nand NAND2_304(II2577,WX1002,WX683);
  nand NAND2_305(II2578,WX1002,II2577);
  nand NAND2_306(II2579,WX683,II2577);
  nand NAND2_307(II2576,II2578,II2579);
  nand NAND2_308(II2584,WX747,II2576);
  nand NAND2_309(II2585,WX747,II2584);
  nand NAND2_310(II2586,II2576,II2584);
  nand NAND2_311(II2575,II2585,II2586);
  nand NAND2_312(II2592,WX811,WX875);
  nand NAND2_313(II2593,WX811,II2592);
  nand NAND2_314(II2594,WX875,II2592);
  nand NAND2_315(II2591,II2593,II2594);
  nand NAND2_316(II2599,II2575,II2591);
  nand NAND2_317(II2600,II2575,II2599);
  nand NAND2_318(II2601,II2591,II2599);
  nand NAND2_319(WX919,II2600,II2601);
  nand NAND2_320(II2608,WX1002,WX685);
  nand NAND2_321(II2609,WX1002,II2608);
  nand NAND2_322(II2610,WX685,II2608);
  nand NAND2_323(II2607,II2609,II2610);
  nand NAND2_324(II2615,WX749,II2607);
  nand NAND2_325(II2616,WX749,II2615);
  nand NAND2_326(II2617,II2607,II2615);
  nand NAND2_327(II2606,II2616,II2617);
  nand NAND2_328(II2623,WX813,WX877);
  nand NAND2_329(II2624,WX813,II2623);
  nand NAND2_330(II2625,WX877,II2623);
  nand NAND2_331(II2622,II2624,II2625);
  nand NAND2_332(II2630,II2606,II2622);
  nand NAND2_333(II2631,II2606,II2630);
  nand NAND2_334(II2632,II2622,II2630);
  nand NAND2_335(WX920,II2631,II2632);
  nand NAND2_336(II2639,WX1002,WX687);
  nand NAND2_337(II2640,WX1002,II2639);
  nand NAND2_338(II2641,WX687,II2639);
  nand NAND2_339(II2638,II2640,II2641);
  nand NAND2_340(II2646,WX751,II2638);
  nand NAND2_341(II2647,WX751,II2646);
  nand NAND2_342(II2648,II2638,II2646);
  nand NAND2_343(II2637,II2647,II2648);
  nand NAND2_344(II2654,WX815,WX879);
  nand NAND2_345(II2655,WX815,II2654);
  nand NAND2_346(II2656,WX879,II2654);
  nand NAND2_347(II2653,II2655,II2656);
  nand NAND2_348(II2661,II2637,II2653);
  nand NAND2_349(II2662,II2637,II2661);
  nand NAND2_350(II2663,II2653,II2661);
  nand NAND2_351(WX921,II2662,II2663);
  nand NAND2_352(II2670,WX1002,WX689);
  nand NAND2_353(II2671,WX1002,II2670);
  nand NAND2_354(II2672,WX689,II2670);
  nand NAND2_355(II2669,II2671,II2672);
  nand NAND2_356(II2677,WX753,II2669);
  nand NAND2_357(II2678,WX753,II2677);
  nand NAND2_358(II2679,II2669,II2677);
  nand NAND2_359(II2668,II2678,II2679);
  nand NAND2_360(II2685,WX817,WX881);
  nand NAND2_361(II2686,WX817,II2685);
  nand NAND2_362(II2687,WX881,II2685);
  nand NAND2_363(II2684,II2686,II2687);
  nand NAND2_364(II2692,II2668,II2684);
  nand NAND2_365(II2693,II2668,II2692);
  nand NAND2_366(II2694,II2684,II2692);
  nand NAND2_367(WX922,II2693,II2694);
  nand NAND2_368(II2701,WX1002,WX691);
  nand NAND2_369(II2702,WX1002,II2701);
  nand NAND2_370(II2703,WX691,II2701);
  nand NAND2_371(II2700,II2702,II2703);
  nand NAND2_372(II2708,WX755,II2700);
  nand NAND2_373(II2709,WX755,II2708);
  nand NAND2_374(II2710,II2700,II2708);
  nand NAND2_375(II2699,II2709,II2710);
  nand NAND2_376(II2716,WX819,WX883);
  nand NAND2_377(II2717,WX819,II2716);
  nand NAND2_378(II2718,WX883,II2716);
  nand NAND2_379(II2715,II2717,II2718);
  nand NAND2_380(II2723,II2699,II2715);
  nand NAND2_381(II2724,II2699,II2723);
  nand NAND2_382(II2725,II2715,II2723);
  nand NAND2_383(WX923,II2724,II2725);
  nand NAND2_384(II2732,WX1002,WX693);
  nand NAND2_385(II2733,WX1002,II2732);
  nand NAND2_386(II2734,WX693,II2732);
  nand NAND2_387(II2731,II2733,II2734);
  nand NAND2_388(II2739,WX757,II2731);
  nand NAND2_389(II2740,WX757,II2739);
  nand NAND2_390(II2741,II2731,II2739);
  nand NAND2_391(II2730,II2740,II2741);
  nand NAND2_392(II2747,WX821,WX885);
  nand NAND2_393(II2748,WX821,II2747);
  nand NAND2_394(II2749,WX885,II2747);
  nand NAND2_395(II2746,II2748,II2749);
  nand NAND2_396(II2754,II2730,II2746);
  nand NAND2_397(II2755,II2730,II2754);
  nand NAND2_398(II2756,II2746,II2754);
  nand NAND2_399(WX924,II2755,II2756);
  nand NAND2_400(II2763,WX1002,WX695);
  nand NAND2_401(II2764,WX1002,II2763);
  nand NAND2_402(II2765,WX695,II2763);
  nand NAND2_403(II2762,II2764,II2765);
  nand NAND2_404(II2770,WX759,II2762);
  nand NAND2_405(II2771,WX759,II2770);
  nand NAND2_406(II2772,II2762,II2770);
  nand NAND2_407(II2761,II2771,II2772);
  nand NAND2_408(II2778,WX823,WX887);
  nand NAND2_409(II2779,WX823,II2778);
  nand NAND2_410(II2780,WX887,II2778);
  nand NAND2_411(II2777,II2779,II2780);
  nand NAND2_412(II2785,II2761,II2777);
  nand NAND2_413(II2786,II2761,II2785);
  nand NAND2_414(II2787,II2777,II2785);
  nand NAND2_415(WX925,II2786,II2787);
  nand NAND2_416(II2794,WX1002,WX697);
  nand NAND2_417(II2795,WX1002,II2794);
  nand NAND2_418(II2796,WX697,II2794);
  nand NAND2_419(II2793,II2795,II2796);
  nand NAND2_420(II2801,WX761,II2793);
  nand NAND2_421(II2802,WX761,II2801);
  nand NAND2_422(II2803,II2793,II2801);
  nand NAND2_423(II2792,II2802,II2803);
  nand NAND2_424(II2809,WX825,WX889);
  nand NAND2_425(II2810,WX825,II2809);
  nand NAND2_426(II2811,WX889,II2809);
  nand NAND2_427(II2808,II2810,II2811);
  nand NAND2_428(II2816,II2792,II2808);
  nand NAND2_429(II2817,II2792,II2816);
  nand NAND2_430(II2818,II2808,II2816);
  nand NAND2_431(WX926,II2817,II2818);
  nand NAND2_432(II2825,WX1002,WX699);
  nand NAND2_433(II2826,WX1002,II2825);
  nand NAND2_434(II2827,WX699,II2825);
  nand NAND2_435(II2824,II2826,II2827);
  nand NAND2_436(II2832,WX763,II2824);
  nand NAND2_437(II2833,WX763,II2832);
  nand NAND2_438(II2834,II2824,II2832);
  nand NAND2_439(II2823,II2833,II2834);
  nand NAND2_440(II2840,WX827,WX891);
  nand NAND2_441(II2841,WX827,II2840);
  nand NAND2_442(II2842,WX891,II2840);
  nand NAND2_443(II2839,II2841,II2842);
  nand NAND2_444(II2847,II2823,II2839);
  nand NAND2_445(II2848,II2823,II2847);
  nand NAND2_446(II2849,II2839,II2847);
  nand NAND2_447(WX927,II2848,II2849);
  nand NAND2_448(II2856,WX1002,WX701);
  nand NAND2_449(II2857,WX1002,II2856);
  nand NAND2_450(II2858,WX701,II2856);
  nand NAND2_451(II2855,II2857,II2858);
  nand NAND2_452(II2863,WX765,II2855);
  nand NAND2_453(II2864,WX765,II2863);
  nand NAND2_454(II2865,II2855,II2863);
  nand NAND2_455(II2854,II2864,II2865);
  nand NAND2_456(II2871,WX829,WX893);
  nand NAND2_457(II2872,WX829,II2871);
  nand NAND2_458(II2873,WX893,II2871);
  nand NAND2_459(II2870,II2872,II2873);
  nand NAND2_460(II2878,II2854,II2870);
  nand NAND2_461(II2879,II2854,II2878);
  nand NAND2_462(II2880,II2870,II2878);
  nand NAND2_463(WX928,II2879,II2880);
  nand NAND2_464(II2887,WX1002,WX703);
  nand NAND2_465(II2888,WX1002,II2887);
  nand NAND2_466(II2889,WX703,II2887);
  nand NAND2_467(II2886,II2888,II2889);
  nand NAND2_468(II2894,WX767,II2886);
  nand NAND2_469(II2895,WX767,II2894);
  nand NAND2_470(II2896,II2886,II2894);
  nand NAND2_471(II2885,II2895,II2896);
  nand NAND2_472(II2902,WX831,WX895);
  nand NAND2_473(II2903,WX831,II2902);
  nand NAND2_474(II2904,WX895,II2902);
  nand NAND2_475(II2901,II2903,II2904);
  nand NAND2_476(II2909,II2885,II2901);
  nand NAND2_477(II2910,II2885,II2909);
  nand NAND2_478(II2911,II2901,II2909);
  nand NAND2_479(WX929,II2910,II2911);
  nand NAND2_480(II2918,WX1002,WX705);
  nand NAND2_481(II2919,WX1002,II2918);
  nand NAND2_482(II2920,WX705,II2918);
  nand NAND2_483(II2917,II2919,II2920);
  nand NAND2_484(II2925,WX769,II2917);
  nand NAND2_485(II2926,WX769,II2925);
  nand NAND2_486(II2927,II2917,II2925);
  nand NAND2_487(II2916,II2926,II2927);
  nand NAND2_488(II2933,WX833,WX897);
  nand NAND2_489(II2934,WX833,II2933);
  nand NAND2_490(II2935,WX897,II2933);
  nand NAND2_491(II2932,II2934,II2935);
  nand NAND2_492(II2940,II2916,II2932);
  nand NAND2_493(II2941,II2916,II2940);
  nand NAND2_494(II2942,II2932,II2940);
  nand NAND2_495(WX930,II2941,II2942);
  nand NAND2_496(II2949,WX1002,WX707);
  nand NAND2_497(II2950,WX1002,II2949);
  nand NAND2_498(II2951,WX707,II2949);
  nand NAND2_499(II2948,II2950,II2951);
  nand NAND2_500(II2956,WX771,II2948);
  nand NAND2_501(II2957,WX771,II2956);
  nand NAND2_502(II2958,II2948,II2956);
  nand NAND2_503(II2947,II2957,II2958);
  nand NAND2_504(II2964,WX835,WX899);
  nand NAND2_505(II2965,WX835,II2964);
  nand NAND2_506(II2966,WX899,II2964);
  nand NAND2_507(II2963,II2965,II2966);
  nand NAND2_508(II2971,II2947,II2963);
  nand NAND2_509(II2972,II2947,II2971);
  nand NAND2_510(II2973,II2963,II2971);
  nand NAND2_511(WX931,II2972,II2973);
  nand NAND2_512(II3052,WX580,WX485);
  nand NAND2_513(II3053,WX580,II3052);
  nand NAND2_514(II3054,WX485,II3052);
  nand NAND2_515(WX1006,II3053,II3054);
  nand NAND2_516(II3065,WX581,WX487);
  nand NAND2_517(II3066,WX581,II3065);
  nand NAND2_518(II3067,WX487,II3065);
  nand NAND2_519(WX1013,II3066,II3067);
  nand NAND2_520(II3078,WX582,WX489);
  nand NAND2_521(II3079,WX582,II3078);
  nand NAND2_522(II3080,WX489,II3078);
  nand NAND2_523(WX1020,II3079,II3080);
  nand NAND2_524(II3091,WX583,WX491);
  nand NAND2_525(II3092,WX583,II3091);
  nand NAND2_526(II3093,WX491,II3091);
  nand NAND2_527(WX1027,II3092,II3093);
  nand NAND2_528(II3104,WX584,WX493);
  nand NAND2_529(II3105,WX584,II3104);
  nand NAND2_530(II3106,WX493,II3104);
  nand NAND2_531(WX1034,II3105,II3106);
  nand NAND2_532(II3117,WX585,WX495);
  nand NAND2_533(II3118,WX585,II3117);
  nand NAND2_534(II3119,WX495,II3117);
  nand NAND2_535(WX1041,II3118,II3119);
  nand NAND2_536(II3130,WX586,WX497);
  nand NAND2_537(II3131,WX586,II3130);
  nand NAND2_538(II3132,WX497,II3130);
  nand NAND2_539(WX1048,II3131,II3132);
  nand NAND2_540(II3143,WX587,WX499);
  nand NAND2_541(II3144,WX587,II3143);
  nand NAND2_542(II3145,WX499,II3143);
  nand NAND2_543(WX1055,II3144,II3145);
  nand NAND2_544(II3156,WX588,WX501);
  nand NAND2_545(II3157,WX588,II3156);
  nand NAND2_546(II3158,WX501,II3156);
  nand NAND2_547(WX1062,II3157,II3158);
  nand NAND2_548(II3169,WX589,WX503);
  nand NAND2_549(II3170,WX589,II3169);
  nand NAND2_550(II3171,WX503,II3169);
  nand NAND2_551(WX1069,II3170,II3171);
  nand NAND2_552(II3182,WX590,WX505);
  nand NAND2_553(II3183,WX590,II3182);
  nand NAND2_554(II3184,WX505,II3182);
  nand NAND2_555(WX1076,II3183,II3184);
  nand NAND2_556(II3195,WX591,WX507);
  nand NAND2_557(II3196,WX591,II3195);
  nand NAND2_558(II3197,WX507,II3195);
  nand NAND2_559(WX1083,II3196,II3197);
  nand NAND2_560(II3208,WX592,WX509);
  nand NAND2_561(II3209,WX592,II3208);
  nand NAND2_562(II3210,WX509,II3208);
  nand NAND2_563(WX1090,II3209,II3210);
  nand NAND2_564(II3221,WX593,WX511);
  nand NAND2_565(II3222,WX593,II3221);
  nand NAND2_566(II3223,WX511,II3221);
  nand NAND2_567(WX1097,II3222,II3223);
  nand NAND2_568(II3234,WX594,WX513);
  nand NAND2_569(II3235,WX594,II3234);
  nand NAND2_570(II3236,WX513,II3234);
  nand NAND2_571(WX1104,II3235,II3236);
  nand NAND2_572(II3247,WX595,WX515);
  nand NAND2_573(II3248,WX595,II3247);
  nand NAND2_574(II3249,WX515,II3247);
  nand NAND2_575(WX1111,II3248,II3249);
  nand NAND2_576(II3260,WX596,WX517);
  nand NAND2_577(II3261,WX596,II3260);
  nand NAND2_578(II3262,WX517,II3260);
  nand NAND2_579(WX1118,II3261,II3262);
  nand NAND2_580(II3273,WX597,WX519);
  nand NAND2_581(II3274,WX597,II3273);
  nand NAND2_582(II3275,WX519,II3273);
  nand NAND2_583(WX1125,II3274,II3275);
  nand NAND2_584(II3286,WX598,WX521);
  nand NAND2_585(II3287,WX598,II3286);
  nand NAND2_586(II3288,WX521,II3286);
  nand NAND2_587(WX1132,II3287,II3288);
  nand NAND2_588(II3299,WX599,WX523);
  nand NAND2_589(II3300,WX599,II3299);
  nand NAND2_590(II3301,WX523,II3299);
  nand NAND2_591(WX1139,II3300,II3301);
  nand NAND2_592(II3312,WX600,WX525);
  nand NAND2_593(II3313,WX600,II3312);
  nand NAND2_594(II3314,WX525,II3312);
  nand NAND2_595(WX1146,II3313,II3314);
  nand NAND2_596(II3325,WX601,WX527);
  nand NAND2_597(II3326,WX601,II3325);
  nand NAND2_598(II3327,WX527,II3325);
  nand NAND2_599(WX1153,II3326,II3327);
  nand NAND2_600(II3338,WX602,WX529);
  nand NAND2_601(II3339,WX602,II3338);
  nand NAND2_602(II3340,WX529,II3338);
  nand NAND2_603(WX1160,II3339,II3340);
  nand NAND2_604(II3351,WX603,WX531);
  nand NAND2_605(II3352,WX603,II3351);
  nand NAND2_606(II3353,WX531,II3351);
  nand NAND2_607(WX1167,II3352,II3353);
  nand NAND2_608(II3364,WX604,WX533);
  nand NAND2_609(II3365,WX604,II3364);
  nand NAND2_610(II3366,WX533,II3364);
  nand NAND2_611(WX1174,II3365,II3366);
  nand NAND2_612(II3377,WX605,WX535);
  nand NAND2_613(II3378,WX605,II3377);
  nand NAND2_614(II3379,WX535,II3377);
  nand NAND2_615(WX1181,II3378,II3379);
  nand NAND2_616(II3390,WX606,WX537);
  nand NAND2_617(II3391,WX606,II3390);
  nand NAND2_618(II3392,WX537,II3390);
  nand NAND2_619(WX1188,II3391,II3392);
  nand NAND2_620(II3403,WX607,WX539);
  nand NAND2_621(II3404,WX607,II3403);
  nand NAND2_622(II3405,WX539,II3403);
  nand NAND2_623(WX1195,II3404,II3405);
  nand NAND2_624(II3416,WX608,WX541);
  nand NAND2_625(II3417,WX608,II3416);
  nand NAND2_626(II3418,WX541,II3416);
  nand NAND2_627(WX1202,II3417,II3418);
  nand NAND2_628(II3429,WX609,WX543);
  nand NAND2_629(II3430,WX609,II3429);
  nand NAND2_630(II3431,WX543,II3429);
  nand NAND2_631(WX1209,II3430,II3431);
  nand NAND2_632(II3442,WX610,WX545);
  nand NAND2_633(II3443,WX610,II3442);
  nand NAND2_634(II3444,WX545,II3442);
  nand NAND2_635(WX1216,II3443,II3444);
  nand NAND2_636(II3455,WX611,WX547);
  nand NAND2_637(II3456,WX611,II3455);
  nand NAND2_638(II3457,WX547,II3455);
  nand NAND2_639(WX1223,II3456,II3457);
  nand NAND2_640(II3470,WX627,CRC_OUT_9_31);
  nand NAND2_641(II3471,WX627,II3470);
  nand NAND2_642(II3472,CRC_OUT_9_31,II3470);
  nand NAND2_643(II3469,II3471,II3472);
  nand NAND2_644(II3477,CRC_OUT_9_15,II3469);
  nand NAND2_645(II3478,CRC_OUT_9_15,II3477);
  nand NAND2_646(II3479,II3469,II3477);
  nand NAND2_647(WX1231,II3478,II3479);
  nand NAND2_648(II3485,WX632,CRC_OUT_9_31);
  nand NAND2_649(II3486,WX632,II3485);
  nand NAND2_650(II3487,CRC_OUT_9_31,II3485);
  nand NAND2_651(II3484,II3486,II3487);
  nand NAND2_652(II3492,CRC_OUT_9_10,II3484);
  nand NAND2_653(II3493,CRC_OUT_9_10,II3492);
  nand NAND2_654(II3494,II3484,II3492);
  nand NAND2_655(WX1232,II3493,II3494);
  nand NAND2_656(II3500,WX639,CRC_OUT_9_31);
  nand NAND2_657(II3501,WX639,II3500);
  nand NAND2_658(II3502,CRC_OUT_9_31,II3500);
  nand NAND2_659(II3499,II3501,II3502);
  nand NAND2_660(II3507,CRC_OUT_9_3,II3499);
  nand NAND2_661(II3508,CRC_OUT_9_3,II3507);
  nand NAND2_662(II3509,II3499,II3507);
  nand NAND2_663(WX1233,II3508,II3509);
  nand NAND2_664(II3514,WX643,CRC_OUT_9_31);
  nand NAND2_665(II3515,WX643,II3514);
  nand NAND2_666(II3516,CRC_OUT_9_31,II3514);
  nand NAND2_667(WX1234,II3515,II3516);
  nand NAND2_668(II3521,WX612,CRC_OUT_9_30);
  nand NAND2_669(II3522,WX612,II3521);
  nand NAND2_670(II3523,CRC_OUT_9_30,II3521);
  nand NAND2_671(WX1235,II3522,II3523);
  nand NAND2_672(II3528,WX613,CRC_OUT_9_29);
  nand NAND2_673(II3529,WX613,II3528);
  nand NAND2_674(II3530,CRC_OUT_9_29,II3528);
  nand NAND2_675(WX1236,II3529,II3530);
  nand NAND2_676(II3535,WX614,CRC_OUT_9_28);
  nand NAND2_677(II3536,WX614,II3535);
  nand NAND2_678(II3537,CRC_OUT_9_28,II3535);
  nand NAND2_679(WX1237,II3536,II3537);
  nand NAND2_680(II3542,WX615,CRC_OUT_9_27);
  nand NAND2_681(II3543,WX615,II3542);
  nand NAND2_682(II3544,CRC_OUT_9_27,II3542);
  nand NAND2_683(WX1238,II3543,II3544);
  nand NAND2_684(II3549,WX616,CRC_OUT_9_26);
  nand NAND2_685(II3550,WX616,II3549);
  nand NAND2_686(II3551,CRC_OUT_9_26,II3549);
  nand NAND2_687(WX1239,II3550,II3551);
  nand NAND2_688(II3556,WX617,CRC_OUT_9_25);
  nand NAND2_689(II3557,WX617,II3556);
  nand NAND2_690(II3558,CRC_OUT_9_25,II3556);
  nand NAND2_691(WX1240,II3557,II3558);
  nand NAND2_692(II3563,WX618,CRC_OUT_9_24);
  nand NAND2_693(II3564,WX618,II3563);
  nand NAND2_694(II3565,CRC_OUT_9_24,II3563);
  nand NAND2_695(WX1241,II3564,II3565);
  nand NAND2_696(II3570,WX619,CRC_OUT_9_23);
  nand NAND2_697(II3571,WX619,II3570);
  nand NAND2_698(II3572,CRC_OUT_9_23,II3570);
  nand NAND2_699(WX1242,II3571,II3572);
  nand NAND2_700(II3577,WX620,CRC_OUT_9_22);
  nand NAND2_701(II3578,WX620,II3577);
  nand NAND2_702(II3579,CRC_OUT_9_22,II3577);
  nand NAND2_703(WX1243,II3578,II3579);
  nand NAND2_704(II3584,WX621,CRC_OUT_9_21);
  nand NAND2_705(II3585,WX621,II3584);
  nand NAND2_706(II3586,CRC_OUT_9_21,II3584);
  nand NAND2_707(WX1244,II3585,II3586);
  nand NAND2_708(II3591,WX622,CRC_OUT_9_20);
  nand NAND2_709(II3592,WX622,II3591);
  nand NAND2_710(II3593,CRC_OUT_9_20,II3591);
  nand NAND2_711(WX1245,II3592,II3593);
  nand NAND2_712(II3598,WX623,CRC_OUT_9_19);
  nand NAND2_713(II3599,WX623,II3598);
  nand NAND2_714(II3600,CRC_OUT_9_19,II3598);
  nand NAND2_715(WX1246,II3599,II3600);
  nand NAND2_716(II3605,WX624,CRC_OUT_9_18);
  nand NAND2_717(II3606,WX624,II3605);
  nand NAND2_718(II3607,CRC_OUT_9_18,II3605);
  nand NAND2_719(WX1247,II3606,II3607);
  nand NAND2_720(II3612,WX625,CRC_OUT_9_17);
  nand NAND2_721(II3613,WX625,II3612);
  nand NAND2_722(II3614,CRC_OUT_9_17,II3612);
  nand NAND2_723(WX1248,II3613,II3614);
  nand NAND2_724(II3619,WX626,CRC_OUT_9_16);
  nand NAND2_725(II3620,WX626,II3619);
  nand NAND2_726(II3621,CRC_OUT_9_16,II3619);
  nand NAND2_727(WX1249,II3620,II3621);
  nand NAND2_728(II3626,WX628,CRC_OUT_9_14);
  nand NAND2_729(II3627,WX628,II3626);
  nand NAND2_730(II3628,CRC_OUT_9_14,II3626);
  nand NAND2_731(WX1250,II3627,II3628);
  nand NAND2_732(II3633,WX629,CRC_OUT_9_13);
  nand NAND2_733(II3634,WX629,II3633);
  nand NAND2_734(II3635,CRC_OUT_9_13,II3633);
  nand NAND2_735(WX1251,II3634,II3635);
  nand NAND2_736(II3640,WX630,CRC_OUT_9_12);
  nand NAND2_737(II3641,WX630,II3640);
  nand NAND2_738(II3642,CRC_OUT_9_12,II3640);
  nand NAND2_739(WX1252,II3641,II3642);
  nand NAND2_740(II3647,WX631,CRC_OUT_9_11);
  nand NAND2_741(II3648,WX631,II3647);
  nand NAND2_742(II3649,CRC_OUT_9_11,II3647);
  nand NAND2_743(WX1253,II3648,II3649);
  nand NAND2_744(II3654,WX633,CRC_OUT_9_9);
  nand NAND2_745(II3655,WX633,II3654);
  nand NAND2_746(II3656,CRC_OUT_9_9,II3654);
  nand NAND2_747(WX1254,II3655,II3656);
  nand NAND2_748(II3661,WX634,CRC_OUT_9_8);
  nand NAND2_749(II3662,WX634,II3661);
  nand NAND2_750(II3663,CRC_OUT_9_8,II3661);
  nand NAND2_751(WX1255,II3662,II3663);
  nand NAND2_752(II3668,WX635,CRC_OUT_9_7);
  nand NAND2_753(II3669,WX635,II3668);
  nand NAND2_754(II3670,CRC_OUT_9_7,II3668);
  nand NAND2_755(WX1256,II3669,II3670);
  nand NAND2_756(II3675,WX636,CRC_OUT_9_6);
  nand NAND2_757(II3676,WX636,II3675);
  nand NAND2_758(II3677,CRC_OUT_9_6,II3675);
  nand NAND2_759(WX1257,II3676,II3677);
  nand NAND2_760(II3682,WX637,CRC_OUT_9_5);
  nand NAND2_761(II3683,WX637,II3682);
  nand NAND2_762(II3684,CRC_OUT_9_5,II3682);
  nand NAND2_763(WX1258,II3683,II3684);
  nand NAND2_764(II3689,WX638,CRC_OUT_9_4);
  nand NAND2_765(II3690,WX638,II3689);
  nand NAND2_766(II3691,CRC_OUT_9_4,II3689);
  nand NAND2_767(WX1259,II3690,II3691);
  nand NAND2_768(II3696,WX640,CRC_OUT_9_2);
  nand NAND2_769(II3697,WX640,II3696);
  nand NAND2_770(II3698,CRC_OUT_9_2,II3696);
  nand NAND2_771(WX1260,II3697,II3698);
  nand NAND2_772(II3703,WX641,CRC_OUT_9_1);
  nand NAND2_773(II3704,WX641,II3703);
  nand NAND2_774(II3705,CRC_OUT_9_1,II3703);
  nand NAND2_775(WX1261,II3704,II3705);
  nand NAND2_776(II3710,WX642,CRC_OUT_9_0);
  nand NAND2_777(II3711,WX642,II3710);
  nand NAND2_778(II3712,CRC_OUT_9_0,II3710);
  nand NAND2_779(WX1262,II3711,II3712);
  nand NAND2_780(II5993,WX2294,WX1938);
  nand NAND2_781(II5994,WX2294,II5993);
  nand NAND2_782(II5995,WX1938,II5993);
  nand NAND2_783(II5992,II5994,II5995);
  nand NAND2_784(II6000,WX2002,II5992);
  nand NAND2_785(II6001,WX2002,II6000);
  nand NAND2_786(II6002,II5992,II6000);
  nand NAND2_787(II5991,II6001,II6002);
  nand NAND2_788(II6008,WX2066,WX2130);
  nand NAND2_789(II6009,WX2066,II6008);
  nand NAND2_790(II6010,WX2130,II6008);
  nand NAND2_791(II6007,II6009,II6010);
  nand NAND2_792(II6015,II5991,II6007);
  nand NAND2_793(II6016,II5991,II6015);
  nand NAND2_794(II6017,II6007,II6015);
  nand NAND2_795(WX2193,II6016,II6017);
  nand NAND2_796(II6024,WX2294,WX1940);
  nand NAND2_797(II6025,WX2294,II6024);
  nand NAND2_798(II6026,WX1940,II6024);
  nand NAND2_799(II6023,II6025,II6026);
  nand NAND2_800(II6031,WX2004,II6023);
  nand NAND2_801(II6032,WX2004,II6031);
  nand NAND2_802(II6033,II6023,II6031);
  nand NAND2_803(II6022,II6032,II6033);
  nand NAND2_804(II6039,WX2068,WX2132);
  nand NAND2_805(II6040,WX2068,II6039);
  nand NAND2_806(II6041,WX2132,II6039);
  nand NAND2_807(II6038,II6040,II6041);
  nand NAND2_808(II6046,II6022,II6038);
  nand NAND2_809(II6047,II6022,II6046);
  nand NAND2_810(II6048,II6038,II6046);
  nand NAND2_811(WX2194,II6047,II6048);
  nand NAND2_812(II6055,WX2294,WX1942);
  nand NAND2_813(II6056,WX2294,II6055);
  nand NAND2_814(II6057,WX1942,II6055);
  nand NAND2_815(II6054,II6056,II6057);
  nand NAND2_816(II6062,WX2006,II6054);
  nand NAND2_817(II6063,WX2006,II6062);
  nand NAND2_818(II6064,II6054,II6062);
  nand NAND2_819(II6053,II6063,II6064);
  nand NAND2_820(II6070,WX2070,WX2134);
  nand NAND2_821(II6071,WX2070,II6070);
  nand NAND2_822(II6072,WX2134,II6070);
  nand NAND2_823(II6069,II6071,II6072);
  nand NAND2_824(II6077,II6053,II6069);
  nand NAND2_825(II6078,II6053,II6077);
  nand NAND2_826(II6079,II6069,II6077);
  nand NAND2_827(WX2195,II6078,II6079);
  nand NAND2_828(II6086,WX2294,WX1944);
  nand NAND2_829(II6087,WX2294,II6086);
  nand NAND2_830(II6088,WX1944,II6086);
  nand NAND2_831(II6085,II6087,II6088);
  nand NAND2_832(II6093,WX2008,II6085);
  nand NAND2_833(II6094,WX2008,II6093);
  nand NAND2_834(II6095,II6085,II6093);
  nand NAND2_835(II6084,II6094,II6095);
  nand NAND2_836(II6101,WX2072,WX2136);
  nand NAND2_837(II6102,WX2072,II6101);
  nand NAND2_838(II6103,WX2136,II6101);
  nand NAND2_839(II6100,II6102,II6103);
  nand NAND2_840(II6108,II6084,II6100);
  nand NAND2_841(II6109,II6084,II6108);
  nand NAND2_842(II6110,II6100,II6108);
  nand NAND2_843(WX2196,II6109,II6110);
  nand NAND2_844(II6117,WX2294,WX1946);
  nand NAND2_845(II6118,WX2294,II6117);
  nand NAND2_846(II6119,WX1946,II6117);
  nand NAND2_847(II6116,II6118,II6119);
  nand NAND2_848(II6124,WX2010,II6116);
  nand NAND2_849(II6125,WX2010,II6124);
  nand NAND2_850(II6126,II6116,II6124);
  nand NAND2_851(II6115,II6125,II6126);
  nand NAND2_852(II6132,WX2074,WX2138);
  nand NAND2_853(II6133,WX2074,II6132);
  nand NAND2_854(II6134,WX2138,II6132);
  nand NAND2_855(II6131,II6133,II6134);
  nand NAND2_856(II6139,II6115,II6131);
  nand NAND2_857(II6140,II6115,II6139);
  nand NAND2_858(II6141,II6131,II6139);
  nand NAND2_859(WX2197,II6140,II6141);
  nand NAND2_860(II6148,WX2294,WX1948);
  nand NAND2_861(II6149,WX2294,II6148);
  nand NAND2_862(II6150,WX1948,II6148);
  nand NAND2_863(II6147,II6149,II6150);
  nand NAND2_864(II6155,WX2012,II6147);
  nand NAND2_865(II6156,WX2012,II6155);
  nand NAND2_866(II6157,II6147,II6155);
  nand NAND2_867(II6146,II6156,II6157);
  nand NAND2_868(II6163,WX2076,WX2140);
  nand NAND2_869(II6164,WX2076,II6163);
  nand NAND2_870(II6165,WX2140,II6163);
  nand NAND2_871(II6162,II6164,II6165);
  nand NAND2_872(II6170,II6146,II6162);
  nand NAND2_873(II6171,II6146,II6170);
  nand NAND2_874(II6172,II6162,II6170);
  nand NAND2_875(WX2198,II6171,II6172);
  nand NAND2_876(II6179,WX2294,WX1950);
  nand NAND2_877(II6180,WX2294,II6179);
  nand NAND2_878(II6181,WX1950,II6179);
  nand NAND2_879(II6178,II6180,II6181);
  nand NAND2_880(II6186,WX2014,II6178);
  nand NAND2_881(II6187,WX2014,II6186);
  nand NAND2_882(II6188,II6178,II6186);
  nand NAND2_883(II6177,II6187,II6188);
  nand NAND2_884(II6194,WX2078,WX2142);
  nand NAND2_885(II6195,WX2078,II6194);
  nand NAND2_886(II6196,WX2142,II6194);
  nand NAND2_887(II6193,II6195,II6196);
  nand NAND2_888(II6201,II6177,II6193);
  nand NAND2_889(II6202,II6177,II6201);
  nand NAND2_890(II6203,II6193,II6201);
  nand NAND2_891(WX2199,II6202,II6203);
  nand NAND2_892(II6210,WX2294,WX1952);
  nand NAND2_893(II6211,WX2294,II6210);
  nand NAND2_894(II6212,WX1952,II6210);
  nand NAND2_895(II6209,II6211,II6212);
  nand NAND2_896(II6217,WX2016,II6209);
  nand NAND2_897(II6218,WX2016,II6217);
  nand NAND2_898(II6219,II6209,II6217);
  nand NAND2_899(II6208,II6218,II6219);
  nand NAND2_900(II6225,WX2080,WX2144);
  nand NAND2_901(II6226,WX2080,II6225);
  nand NAND2_902(II6227,WX2144,II6225);
  nand NAND2_903(II6224,II6226,II6227);
  nand NAND2_904(II6232,II6208,II6224);
  nand NAND2_905(II6233,II6208,II6232);
  nand NAND2_906(II6234,II6224,II6232);
  nand NAND2_907(WX2200,II6233,II6234);
  nand NAND2_908(II6241,WX2294,WX1954);
  nand NAND2_909(II6242,WX2294,II6241);
  nand NAND2_910(II6243,WX1954,II6241);
  nand NAND2_911(II6240,II6242,II6243);
  nand NAND2_912(II6248,WX2018,II6240);
  nand NAND2_913(II6249,WX2018,II6248);
  nand NAND2_914(II6250,II6240,II6248);
  nand NAND2_915(II6239,II6249,II6250);
  nand NAND2_916(II6256,WX2082,WX2146);
  nand NAND2_917(II6257,WX2082,II6256);
  nand NAND2_918(II6258,WX2146,II6256);
  nand NAND2_919(II6255,II6257,II6258);
  nand NAND2_920(II6263,II6239,II6255);
  nand NAND2_921(II6264,II6239,II6263);
  nand NAND2_922(II6265,II6255,II6263);
  nand NAND2_923(WX2201,II6264,II6265);
  nand NAND2_924(II6272,WX2294,WX1956);
  nand NAND2_925(II6273,WX2294,II6272);
  nand NAND2_926(II6274,WX1956,II6272);
  nand NAND2_927(II6271,II6273,II6274);
  nand NAND2_928(II6279,WX2020,II6271);
  nand NAND2_929(II6280,WX2020,II6279);
  nand NAND2_930(II6281,II6271,II6279);
  nand NAND2_931(II6270,II6280,II6281);
  nand NAND2_932(II6287,WX2084,WX2148);
  nand NAND2_933(II6288,WX2084,II6287);
  nand NAND2_934(II6289,WX2148,II6287);
  nand NAND2_935(II6286,II6288,II6289);
  nand NAND2_936(II6294,II6270,II6286);
  nand NAND2_937(II6295,II6270,II6294);
  nand NAND2_938(II6296,II6286,II6294);
  nand NAND2_939(WX2202,II6295,II6296);
  nand NAND2_940(II6303,WX2294,WX1958);
  nand NAND2_941(II6304,WX2294,II6303);
  nand NAND2_942(II6305,WX1958,II6303);
  nand NAND2_943(II6302,II6304,II6305);
  nand NAND2_944(II6310,WX2022,II6302);
  nand NAND2_945(II6311,WX2022,II6310);
  nand NAND2_946(II6312,II6302,II6310);
  nand NAND2_947(II6301,II6311,II6312);
  nand NAND2_948(II6318,WX2086,WX2150);
  nand NAND2_949(II6319,WX2086,II6318);
  nand NAND2_950(II6320,WX2150,II6318);
  nand NAND2_951(II6317,II6319,II6320);
  nand NAND2_952(II6325,II6301,II6317);
  nand NAND2_953(II6326,II6301,II6325);
  nand NAND2_954(II6327,II6317,II6325);
  nand NAND2_955(WX2203,II6326,II6327);
  nand NAND2_956(II6334,WX2294,WX1960);
  nand NAND2_957(II6335,WX2294,II6334);
  nand NAND2_958(II6336,WX1960,II6334);
  nand NAND2_959(II6333,II6335,II6336);
  nand NAND2_960(II6341,WX2024,II6333);
  nand NAND2_961(II6342,WX2024,II6341);
  nand NAND2_962(II6343,II6333,II6341);
  nand NAND2_963(II6332,II6342,II6343);
  nand NAND2_964(II6349,WX2088,WX2152);
  nand NAND2_965(II6350,WX2088,II6349);
  nand NAND2_966(II6351,WX2152,II6349);
  nand NAND2_967(II6348,II6350,II6351);
  nand NAND2_968(II6356,II6332,II6348);
  nand NAND2_969(II6357,II6332,II6356);
  nand NAND2_970(II6358,II6348,II6356);
  nand NAND2_971(WX2204,II6357,II6358);
  nand NAND2_972(II6365,WX2294,WX1962);
  nand NAND2_973(II6366,WX2294,II6365);
  nand NAND2_974(II6367,WX1962,II6365);
  nand NAND2_975(II6364,II6366,II6367);
  nand NAND2_976(II6372,WX2026,II6364);
  nand NAND2_977(II6373,WX2026,II6372);
  nand NAND2_978(II6374,II6364,II6372);
  nand NAND2_979(II6363,II6373,II6374);
  nand NAND2_980(II6380,WX2090,WX2154);
  nand NAND2_981(II6381,WX2090,II6380);
  nand NAND2_982(II6382,WX2154,II6380);
  nand NAND2_983(II6379,II6381,II6382);
  nand NAND2_984(II6387,II6363,II6379);
  nand NAND2_985(II6388,II6363,II6387);
  nand NAND2_986(II6389,II6379,II6387);
  nand NAND2_987(WX2205,II6388,II6389);
  nand NAND2_988(II6396,WX2294,WX1964);
  nand NAND2_989(II6397,WX2294,II6396);
  nand NAND2_990(II6398,WX1964,II6396);
  nand NAND2_991(II6395,II6397,II6398);
  nand NAND2_992(II6403,WX2028,II6395);
  nand NAND2_993(II6404,WX2028,II6403);
  nand NAND2_994(II6405,II6395,II6403);
  nand NAND2_995(II6394,II6404,II6405);
  nand NAND2_996(II6411,WX2092,WX2156);
  nand NAND2_997(II6412,WX2092,II6411);
  nand NAND2_998(II6413,WX2156,II6411);
  nand NAND2_999(II6410,II6412,II6413);
  nand NAND2_1000(II6418,II6394,II6410);
  nand NAND2_1001(II6419,II6394,II6418);
  nand NAND2_1002(II6420,II6410,II6418);
  nand NAND2_1003(WX2206,II6419,II6420);
  nand NAND2_1004(II6427,WX2294,WX1966);
  nand NAND2_1005(II6428,WX2294,II6427);
  nand NAND2_1006(II6429,WX1966,II6427);
  nand NAND2_1007(II6426,II6428,II6429);
  nand NAND2_1008(II6434,WX2030,II6426);
  nand NAND2_1009(II6435,WX2030,II6434);
  nand NAND2_1010(II6436,II6426,II6434);
  nand NAND2_1011(II6425,II6435,II6436);
  nand NAND2_1012(II6442,WX2094,WX2158);
  nand NAND2_1013(II6443,WX2094,II6442);
  nand NAND2_1014(II6444,WX2158,II6442);
  nand NAND2_1015(II6441,II6443,II6444);
  nand NAND2_1016(II6449,II6425,II6441);
  nand NAND2_1017(II6450,II6425,II6449);
  nand NAND2_1018(II6451,II6441,II6449);
  nand NAND2_1019(WX2207,II6450,II6451);
  nand NAND2_1020(II6458,WX2294,WX1968);
  nand NAND2_1021(II6459,WX2294,II6458);
  nand NAND2_1022(II6460,WX1968,II6458);
  nand NAND2_1023(II6457,II6459,II6460);
  nand NAND2_1024(II6465,WX2032,II6457);
  nand NAND2_1025(II6466,WX2032,II6465);
  nand NAND2_1026(II6467,II6457,II6465);
  nand NAND2_1027(II6456,II6466,II6467);
  nand NAND2_1028(II6473,WX2096,WX2160);
  nand NAND2_1029(II6474,WX2096,II6473);
  nand NAND2_1030(II6475,WX2160,II6473);
  nand NAND2_1031(II6472,II6474,II6475);
  nand NAND2_1032(II6480,II6456,II6472);
  nand NAND2_1033(II6481,II6456,II6480);
  nand NAND2_1034(II6482,II6472,II6480);
  nand NAND2_1035(WX2208,II6481,II6482);
  nand NAND2_1036(II6489,WX2295,WX1970);
  nand NAND2_1037(II6490,WX2295,II6489);
  nand NAND2_1038(II6491,WX1970,II6489);
  nand NAND2_1039(II6488,II6490,II6491);
  nand NAND2_1040(II6496,WX2034,II6488);
  nand NAND2_1041(II6497,WX2034,II6496);
  nand NAND2_1042(II6498,II6488,II6496);
  nand NAND2_1043(II6487,II6497,II6498);
  nand NAND2_1044(II6504,WX2098,WX2162);
  nand NAND2_1045(II6505,WX2098,II6504);
  nand NAND2_1046(II6506,WX2162,II6504);
  nand NAND2_1047(II6503,II6505,II6506);
  nand NAND2_1048(II6511,II6487,II6503);
  nand NAND2_1049(II6512,II6487,II6511);
  nand NAND2_1050(II6513,II6503,II6511);
  nand NAND2_1051(WX2209,II6512,II6513);
  nand NAND2_1052(II6520,WX2295,WX1972);
  nand NAND2_1053(II6521,WX2295,II6520);
  nand NAND2_1054(II6522,WX1972,II6520);
  nand NAND2_1055(II6519,II6521,II6522);
  nand NAND2_1056(II6527,WX2036,II6519);
  nand NAND2_1057(II6528,WX2036,II6527);
  nand NAND2_1058(II6529,II6519,II6527);
  nand NAND2_1059(II6518,II6528,II6529);
  nand NAND2_1060(II6535,WX2100,WX2164);
  nand NAND2_1061(II6536,WX2100,II6535);
  nand NAND2_1062(II6537,WX2164,II6535);
  nand NAND2_1063(II6534,II6536,II6537);
  nand NAND2_1064(II6542,II6518,II6534);
  nand NAND2_1065(II6543,II6518,II6542);
  nand NAND2_1066(II6544,II6534,II6542);
  nand NAND2_1067(WX2210,II6543,II6544);
  nand NAND2_1068(II6551,WX2295,WX1974);
  nand NAND2_1069(II6552,WX2295,II6551);
  nand NAND2_1070(II6553,WX1974,II6551);
  nand NAND2_1071(II6550,II6552,II6553);
  nand NAND2_1072(II6558,WX2038,II6550);
  nand NAND2_1073(II6559,WX2038,II6558);
  nand NAND2_1074(II6560,II6550,II6558);
  nand NAND2_1075(II6549,II6559,II6560);
  nand NAND2_1076(II6566,WX2102,WX2166);
  nand NAND2_1077(II6567,WX2102,II6566);
  nand NAND2_1078(II6568,WX2166,II6566);
  nand NAND2_1079(II6565,II6567,II6568);
  nand NAND2_1080(II6573,II6549,II6565);
  nand NAND2_1081(II6574,II6549,II6573);
  nand NAND2_1082(II6575,II6565,II6573);
  nand NAND2_1083(WX2211,II6574,II6575);
  nand NAND2_1084(II6582,WX2295,WX1976);
  nand NAND2_1085(II6583,WX2295,II6582);
  nand NAND2_1086(II6584,WX1976,II6582);
  nand NAND2_1087(II6581,II6583,II6584);
  nand NAND2_1088(II6589,WX2040,II6581);
  nand NAND2_1089(II6590,WX2040,II6589);
  nand NAND2_1090(II6591,II6581,II6589);
  nand NAND2_1091(II6580,II6590,II6591);
  nand NAND2_1092(II6597,WX2104,WX2168);
  nand NAND2_1093(II6598,WX2104,II6597);
  nand NAND2_1094(II6599,WX2168,II6597);
  nand NAND2_1095(II6596,II6598,II6599);
  nand NAND2_1096(II6604,II6580,II6596);
  nand NAND2_1097(II6605,II6580,II6604);
  nand NAND2_1098(II6606,II6596,II6604);
  nand NAND2_1099(WX2212,II6605,II6606);
  nand NAND2_1100(II6613,WX2295,WX1978);
  nand NAND2_1101(II6614,WX2295,II6613);
  nand NAND2_1102(II6615,WX1978,II6613);
  nand NAND2_1103(II6612,II6614,II6615);
  nand NAND2_1104(II6620,WX2042,II6612);
  nand NAND2_1105(II6621,WX2042,II6620);
  nand NAND2_1106(II6622,II6612,II6620);
  nand NAND2_1107(II6611,II6621,II6622);
  nand NAND2_1108(II6628,WX2106,WX2170);
  nand NAND2_1109(II6629,WX2106,II6628);
  nand NAND2_1110(II6630,WX2170,II6628);
  nand NAND2_1111(II6627,II6629,II6630);
  nand NAND2_1112(II6635,II6611,II6627);
  nand NAND2_1113(II6636,II6611,II6635);
  nand NAND2_1114(II6637,II6627,II6635);
  nand NAND2_1115(WX2213,II6636,II6637);
  nand NAND2_1116(II6644,WX2295,WX1980);
  nand NAND2_1117(II6645,WX2295,II6644);
  nand NAND2_1118(II6646,WX1980,II6644);
  nand NAND2_1119(II6643,II6645,II6646);
  nand NAND2_1120(II6651,WX2044,II6643);
  nand NAND2_1121(II6652,WX2044,II6651);
  nand NAND2_1122(II6653,II6643,II6651);
  nand NAND2_1123(II6642,II6652,II6653);
  nand NAND2_1124(II6659,WX2108,WX2172);
  nand NAND2_1125(II6660,WX2108,II6659);
  nand NAND2_1126(II6661,WX2172,II6659);
  nand NAND2_1127(II6658,II6660,II6661);
  nand NAND2_1128(II6666,II6642,II6658);
  nand NAND2_1129(II6667,II6642,II6666);
  nand NAND2_1130(II6668,II6658,II6666);
  nand NAND2_1131(WX2214,II6667,II6668);
  nand NAND2_1132(II6675,WX2295,WX1982);
  nand NAND2_1133(II6676,WX2295,II6675);
  nand NAND2_1134(II6677,WX1982,II6675);
  nand NAND2_1135(II6674,II6676,II6677);
  nand NAND2_1136(II6682,WX2046,II6674);
  nand NAND2_1137(II6683,WX2046,II6682);
  nand NAND2_1138(II6684,II6674,II6682);
  nand NAND2_1139(II6673,II6683,II6684);
  nand NAND2_1140(II6690,WX2110,WX2174);
  nand NAND2_1141(II6691,WX2110,II6690);
  nand NAND2_1142(II6692,WX2174,II6690);
  nand NAND2_1143(II6689,II6691,II6692);
  nand NAND2_1144(II6697,II6673,II6689);
  nand NAND2_1145(II6698,II6673,II6697);
  nand NAND2_1146(II6699,II6689,II6697);
  nand NAND2_1147(WX2215,II6698,II6699);
  nand NAND2_1148(II6706,WX2295,WX1984);
  nand NAND2_1149(II6707,WX2295,II6706);
  nand NAND2_1150(II6708,WX1984,II6706);
  nand NAND2_1151(II6705,II6707,II6708);
  nand NAND2_1152(II6713,WX2048,II6705);
  nand NAND2_1153(II6714,WX2048,II6713);
  nand NAND2_1154(II6715,II6705,II6713);
  nand NAND2_1155(II6704,II6714,II6715);
  nand NAND2_1156(II6721,WX2112,WX2176);
  nand NAND2_1157(II6722,WX2112,II6721);
  nand NAND2_1158(II6723,WX2176,II6721);
  nand NAND2_1159(II6720,II6722,II6723);
  nand NAND2_1160(II6728,II6704,II6720);
  nand NAND2_1161(II6729,II6704,II6728);
  nand NAND2_1162(II6730,II6720,II6728);
  nand NAND2_1163(WX2216,II6729,II6730);
  nand NAND2_1164(II6737,WX2295,WX1986);
  nand NAND2_1165(II6738,WX2295,II6737);
  nand NAND2_1166(II6739,WX1986,II6737);
  nand NAND2_1167(II6736,II6738,II6739);
  nand NAND2_1168(II6744,WX2050,II6736);
  nand NAND2_1169(II6745,WX2050,II6744);
  nand NAND2_1170(II6746,II6736,II6744);
  nand NAND2_1171(II6735,II6745,II6746);
  nand NAND2_1172(II6752,WX2114,WX2178);
  nand NAND2_1173(II6753,WX2114,II6752);
  nand NAND2_1174(II6754,WX2178,II6752);
  nand NAND2_1175(II6751,II6753,II6754);
  nand NAND2_1176(II6759,II6735,II6751);
  nand NAND2_1177(II6760,II6735,II6759);
  nand NAND2_1178(II6761,II6751,II6759);
  nand NAND2_1179(WX2217,II6760,II6761);
  nand NAND2_1180(II6768,WX2295,WX1988);
  nand NAND2_1181(II6769,WX2295,II6768);
  nand NAND2_1182(II6770,WX1988,II6768);
  nand NAND2_1183(II6767,II6769,II6770);
  nand NAND2_1184(II6775,WX2052,II6767);
  nand NAND2_1185(II6776,WX2052,II6775);
  nand NAND2_1186(II6777,II6767,II6775);
  nand NAND2_1187(II6766,II6776,II6777);
  nand NAND2_1188(II6783,WX2116,WX2180);
  nand NAND2_1189(II6784,WX2116,II6783);
  nand NAND2_1190(II6785,WX2180,II6783);
  nand NAND2_1191(II6782,II6784,II6785);
  nand NAND2_1192(II6790,II6766,II6782);
  nand NAND2_1193(II6791,II6766,II6790);
  nand NAND2_1194(II6792,II6782,II6790);
  nand NAND2_1195(WX2218,II6791,II6792);
  nand NAND2_1196(II6799,WX2295,WX1990);
  nand NAND2_1197(II6800,WX2295,II6799);
  nand NAND2_1198(II6801,WX1990,II6799);
  nand NAND2_1199(II6798,II6800,II6801);
  nand NAND2_1200(II6806,WX2054,II6798);
  nand NAND2_1201(II6807,WX2054,II6806);
  nand NAND2_1202(II6808,II6798,II6806);
  nand NAND2_1203(II6797,II6807,II6808);
  nand NAND2_1204(II6814,WX2118,WX2182);
  nand NAND2_1205(II6815,WX2118,II6814);
  nand NAND2_1206(II6816,WX2182,II6814);
  nand NAND2_1207(II6813,II6815,II6816);
  nand NAND2_1208(II6821,II6797,II6813);
  nand NAND2_1209(II6822,II6797,II6821);
  nand NAND2_1210(II6823,II6813,II6821);
  nand NAND2_1211(WX2219,II6822,II6823);
  nand NAND2_1212(II6830,WX2295,WX1992);
  nand NAND2_1213(II6831,WX2295,II6830);
  nand NAND2_1214(II6832,WX1992,II6830);
  nand NAND2_1215(II6829,II6831,II6832);
  nand NAND2_1216(II6837,WX2056,II6829);
  nand NAND2_1217(II6838,WX2056,II6837);
  nand NAND2_1218(II6839,II6829,II6837);
  nand NAND2_1219(II6828,II6838,II6839);
  nand NAND2_1220(II6845,WX2120,WX2184);
  nand NAND2_1221(II6846,WX2120,II6845);
  nand NAND2_1222(II6847,WX2184,II6845);
  nand NAND2_1223(II6844,II6846,II6847);
  nand NAND2_1224(II6852,II6828,II6844);
  nand NAND2_1225(II6853,II6828,II6852);
  nand NAND2_1226(II6854,II6844,II6852);
  nand NAND2_1227(WX2220,II6853,II6854);
  nand NAND2_1228(II6861,WX2295,WX1994);
  nand NAND2_1229(II6862,WX2295,II6861);
  nand NAND2_1230(II6863,WX1994,II6861);
  nand NAND2_1231(II6860,II6862,II6863);
  nand NAND2_1232(II6868,WX2058,II6860);
  nand NAND2_1233(II6869,WX2058,II6868);
  nand NAND2_1234(II6870,II6860,II6868);
  nand NAND2_1235(II6859,II6869,II6870);
  nand NAND2_1236(II6876,WX2122,WX2186);
  nand NAND2_1237(II6877,WX2122,II6876);
  nand NAND2_1238(II6878,WX2186,II6876);
  nand NAND2_1239(II6875,II6877,II6878);
  nand NAND2_1240(II6883,II6859,II6875);
  nand NAND2_1241(II6884,II6859,II6883);
  nand NAND2_1242(II6885,II6875,II6883);
  nand NAND2_1243(WX2221,II6884,II6885);
  nand NAND2_1244(II6892,WX2295,WX1996);
  nand NAND2_1245(II6893,WX2295,II6892);
  nand NAND2_1246(II6894,WX1996,II6892);
  nand NAND2_1247(II6891,II6893,II6894);
  nand NAND2_1248(II6899,WX2060,II6891);
  nand NAND2_1249(II6900,WX2060,II6899);
  nand NAND2_1250(II6901,II6891,II6899);
  nand NAND2_1251(II6890,II6900,II6901);
  nand NAND2_1252(II6907,WX2124,WX2188);
  nand NAND2_1253(II6908,WX2124,II6907);
  nand NAND2_1254(II6909,WX2188,II6907);
  nand NAND2_1255(II6906,II6908,II6909);
  nand NAND2_1256(II6914,II6890,II6906);
  nand NAND2_1257(II6915,II6890,II6914);
  nand NAND2_1258(II6916,II6906,II6914);
  nand NAND2_1259(WX2222,II6915,II6916);
  nand NAND2_1260(II6923,WX2295,WX1998);
  nand NAND2_1261(II6924,WX2295,II6923);
  nand NAND2_1262(II6925,WX1998,II6923);
  nand NAND2_1263(II6922,II6924,II6925);
  nand NAND2_1264(II6930,WX2062,II6922);
  nand NAND2_1265(II6931,WX2062,II6930);
  nand NAND2_1266(II6932,II6922,II6930);
  nand NAND2_1267(II6921,II6931,II6932);
  nand NAND2_1268(II6938,WX2126,WX2190);
  nand NAND2_1269(II6939,WX2126,II6938);
  nand NAND2_1270(II6940,WX2190,II6938);
  nand NAND2_1271(II6937,II6939,II6940);
  nand NAND2_1272(II6945,II6921,II6937);
  nand NAND2_1273(II6946,II6921,II6945);
  nand NAND2_1274(II6947,II6937,II6945);
  nand NAND2_1275(WX2223,II6946,II6947);
  nand NAND2_1276(II6954,WX2295,WX2000);
  nand NAND2_1277(II6955,WX2295,II6954);
  nand NAND2_1278(II6956,WX2000,II6954);
  nand NAND2_1279(II6953,II6955,II6956);
  nand NAND2_1280(II6961,WX2064,II6953);
  nand NAND2_1281(II6962,WX2064,II6961);
  nand NAND2_1282(II6963,II6953,II6961);
  nand NAND2_1283(II6952,II6962,II6963);
  nand NAND2_1284(II6969,WX2128,WX2192);
  nand NAND2_1285(II6970,WX2128,II6969);
  nand NAND2_1286(II6971,WX2192,II6969);
  nand NAND2_1287(II6968,II6970,II6971);
  nand NAND2_1288(II6976,II6952,II6968);
  nand NAND2_1289(II6977,II6952,II6976);
  nand NAND2_1290(II6978,II6968,II6976);
  nand NAND2_1291(WX2224,II6977,II6978);
  nand NAND2_1292(II7057,WX1873,WX1778);
  nand NAND2_1293(II7058,WX1873,II7057);
  nand NAND2_1294(II7059,WX1778,II7057);
  nand NAND2_1295(WX2299,II7058,II7059);
  nand NAND2_1296(II7070,WX1874,WX1780);
  nand NAND2_1297(II7071,WX1874,II7070);
  nand NAND2_1298(II7072,WX1780,II7070);
  nand NAND2_1299(WX2306,II7071,II7072);
  nand NAND2_1300(II7083,WX1875,WX1782);
  nand NAND2_1301(II7084,WX1875,II7083);
  nand NAND2_1302(II7085,WX1782,II7083);
  nand NAND2_1303(WX2313,II7084,II7085);
  nand NAND2_1304(II7096,WX1876,WX1784);
  nand NAND2_1305(II7097,WX1876,II7096);
  nand NAND2_1306(II7098,WX1784,II7096);
  nand NAND2_1307(WX2320,II7097,II7098);
  nand NAND2_1308(II7109,WX1877,WX1786);
  nand NAND2_1309(II7110,WX1877,II7109);
  nand NAND2_1310(II7111,WX1786,II7109);
  nand NAND2_1311(WX2327,II7110,II7111);
  nand NAND2_1312(II7122,WX1878,WX1788);
  nand NAND2_1313(II7123,WX1878,II7122);
  nand NAND2_1314(II7124,WX1788,II7122);
  nand NAND2_1315(WX2334,II7123,II7124);
  nand NAND2_1316(II7135,WX1879,WX1790);
  nand NAND2_1317(II7136,WX1879,II7135);
  nand NAND2_1318(II7137,WX1790,II7135);
  nand NAND2_1319(WX2341,II7136,II7137);
  nand NAND2_1320(II7148,WX1880,WX1792);
  nand NAND2_1321(II7149,WX1880,II7148);
  nand NAND2_1322(II7150,WX1792,II7148);
  nand NAND2_1323(WX2348,II7149,II7150);
  nand NAND2_1324(II7161,WX1881,WX1794);
  nand NAND2_1325(II7162,WX1881,II7161);
  nand NAND2_1326(II7163,WX1794,II7161);
  nand NAND2_1327(WX2355,II7162,II7163);
  nand NAND2_1328(II7174,WX1882,WX1796);
  nand NAND2_1329(II7175,WX1882,II7174);
  nand NAND2_1330(II7176,WX1796,II7174);
  nand NAND2_1331(WX2362,II7175,II7176);
  nand NAND2_1332(II7187,WX1883,WX1798);
  nand NAND2_1333(II7188,WX1883,II7187);
  nand NAND2_1334(II7189,WX1798,II7187);
  nand NAND2_1335(WX2369,II7188,II7189);
  nand NAND2_1336(II7200,WX1884,WX1800);
  nand NAND2_1337(II7201,WX1884,II7200);
  nand NAND2_1338(II7202,WX1800,II7200);
  nand NAND2_1339(WX2376,II7201,II7202);
  nand NAND2_1340(II7213,WX1885,WX1802);
  nand NAND2_1341(II7214,WX1885,II7213);
  nand NAND2_1342(II7215,WX1802,II7213);
  nand NAND2_1343(WX2383,II7214,II7215);
  nand NAND2_1344(II7226,WX1886,WX1804);
  nand NAND2_1345(II7227,WX1886,II7226);
  nand NAND2_1346(II7228,WX1804,II7226);
  nand NAND2_1347(WX2390,II7227,II7228);
  nand NAND2_1348(II7239,WX1887,WX1806);
  nand NAND2_1349(II7240,WX1887,II7239);
  nand NAND2_1350(II7241,WX1806,II7239);
  nand NAND2_1351(WX2397,II7240,II7241);
  nand NAND2_1352(II7252,WX1888,WX1808);
  nand NAND2_1353(II7253,WX1888,II7252);
  nand NAND2_1354(II7254,WX1808,II7252);
  nand NAND2_1355(WX2404,II7253,II7254);
  nand NAND2_1356(II7265,WX1889,WX1810);
  nand NAND2_1357(II7266,WX1889,II7265);
  nand NAND2_1358(II7267,WX1810,II7265);
  nand NAND2_1359(WX2411,II7266,II7267);
  nand NAND2_1360(II7278,WX1890,WX1812);
  nand NAND2_1361(II7279,WX1890,II7278);
  nand NAND2_1362(II7280,WX1812,II7278);
  nand NAND2_1363(WX2418,II7279,II7280);
  nand NAND2_1364(II7291,WX1891,WX1814);
  nand NAND2_1365(II7292,WX1891,II7291);
  nand NAND2_1366(II7293,WX1814,II7291);
  nand NAND2_1367(WX2425,II7292,II7293);
  nand NAND2_1368(II7304,WX1892,WX1816);
  nand NAND2_1369(II7305,WX1892,II7304);
  nand NAND2_1370(II7306,WX1816,II7304);
  nand NAND2_1371(WX2432,II7305,II7306);
  nand NAND2_1372(II7317,WX1893,WX1818);
  nand NAND2_1373(II7318,WX1893,II7317);
  nand NAND2_1374(II7319,WX1818,II7317);
  nand NAND2_1375(WX2439,II7318,II7319);
  nand NAND2_1376(II7330,WX1894,WX1820);
  nand NAND2_1377(II7331,WX1894,II7330);
  nand NAND2_1378(II7332,WX1820,II7330);
  nand NAND2_1379(WX2446,II7331,II7332);
  nand NAND2_1380(II7343,WX1895,WX1822);
  nand NAND2_1381(II7344,WX1895,II7343);
  nand NAND2_1382(II7345,WX1822,II7343);
  nand NAND2_1383(WX2453,II7344,II7345);
  nand NAND2_1384(II7356,WX1896,WX1824);
  nand NAND2_1385(II7357,WX1896,II7356);
  nand NAND2_1386(II7358,WX1824,II7356);
  nand NAND2_1387(WX2460,II7357,II7358);
  nand NAND2_1388(II7369,WX1897,WX1826);
  nand NAND2_1389(II7370,WX1897,II7369);
  nand NAND2_1390(II7371,WX1826,II7369);
  nand NAND2_1391(WX2467,II7370,II7371);
  nand NAND2_1392(II7382,WX1898,WX1828);
  nand NAND2_1393(II7383,WX1898,II7382);
  nand NAND2_1394(II7384,WX1828,II7382);
  nand NAND2_1395(WX2474,II7383,II7384);
  nand NAND2_1396(II7395,WX1899,WX1830);
  nand NAND2_1397(II7396,WX1899,II7395);
  nand NAND2_1398(II7397,WX1830,II7395);
  nand NAND2_1399(WX2481,II7396,II7397);
  nand NAND2_1400(II7408,WX1900,WX1832);
  nand NAND2_1401(II7409,WX1900,II7408);
  nand NAND2_1402(II7410,WX1832,II7408);
  nand NAND2_1403(WX2488,II7409,II7410);
  nand NAND2_1404(II7421,WX1901,WX1834);
  nand NAND2_1405(II7422,WX1901,II7421);
  nand NAND2_1406(II7423,WX1834,II7421);
  nand NAND2_1407(WX2495,II7422,II7423);
  nand NAND2_1408(II7434,WX1902,WX1836);
  nand NAND2_1409(II7435,WX1902,II7434);
  nand NAND2_1410(II7436,WX1836,II7434);
  nand NAND2_1411(WX2502,II7435,II7436);
  nand NAND2_1412(II7447,WX1903,WX1838);
  nand NAND2_1413(II7448,WX1903,II7447);
  nand NAND2_1414(II7449,WX1838,II7447);
  nand NAND2_1415(WX2509,II7448,II7449);
  nand NAND2_1416(II7460,WX1904,WX1840);
  nand NAND2_1417(II7461,WX1904,II7460);
  nand NAND2_1418(II7462,WX1840,II7460);
  nand NAND2_1419(WX2516,II7461,II7462);
  nand NAND2_1420(II7475,WX1920,CRC_OUT_8_31);
  nand NAND2_1421(II7476,WX1920,II7475);
  nand NAND2_1422(II7477,CRC_OUT_8_31,II7475);
  nand NAND2_1423(II7474,II7476,II7477);
  nand NAND2_1424(II7482,CRC_OUT_8_15,II7474);
  nand NAND2_1425(II7483,CRC_OUT_8_15,II7482);
  nand NAND2_1426(II7484,II7474,II7482);
  nand NAND2_1427(WX2524,II7483,II7484);
  nand NAND2_1428(II7490,WX1925,CRC_OUT_8_31);
  nand NAND2_1429(II7491,WX1925,II7490);
  nand NAND2_1430(II7492,CRC_OUT_8_31,II7490);
  nand NAND2_1431(II7489,II7491,II7492);
  nand NAND2_1432(II7497,CRC_OUT_8_10,II7489);
  nand NAND2_1433(II7498,CRC_OUT_8_10,II7497);
  nand NAND2_1434(II7499,II7489,II7497);
  nand NAND2_1435(WX2525,II7498,II7499);
  nand NAND2_1436(II7505,WX1932,CRC_OUT_8_31);
  nand NAND2_1437(II7506,WX1932,II7505);
  nand NAND2_1438(II7507,CRC_OUT_8_31,II7505);
  nand NAND2_1439(II7504,II7506,II7507);
  nand NAND2_1440(II7512,CRC_OUT_8_3,II7504);
  nand NAND2_1441(II7513,CRC_OUT_8_3,II7512);
  nand NAND2_1442(II7514,II7504,II7512);
  nand NAND2_1443(WX2526,II7513,II7514);
  nand NAND2_1444(II7519,WX1936,CRC_OUT_8_31);
  nand NAND2_1445(II7520,WX1936,II7519);
  nand NAND2_1446(II7521,CRC_OUT_8_31,II7519);
  nand NAND2_1447(WX2527,II7520,II7521);
  nand NAND2_1448(II7526,WX1905,CRC_OUT_8_30);
  nand NAND2_1449(II7527,WX1905,II7526);
  nand NAND2_1450(II7528,CRC_OUT_8_30,II7526);
  nand NAND2_1451(WX2528,II7527,II7528);
  nand NAND2_1452(II7533,WX1906,CRC_OUT_8_29);
  nand NAND2_1453(II7534,WX1906,II7533);
  nand NAND2_1454(II7535,CRC_OUT_8_29,II7533);
  nand NAND2_1455(WX2529,II7534,II7535);
  nand NAND2_1456(II7540,WX1907,CRC_OUT_8_28);
  nand NAND2_1457(II7541,WX1907,II7540);
  nand NAND2_1458(II7542,CRC_OUT_8_28,II7540);
  nand NAND2_1459(WX2530,II7541,II7542);
  nand NAND2_1460(II7547,WX1908,CRC_OUT_8_27);
  nand NAND2_1461(II7548,WX1908,II7547);
  nand NAND2_1462(II7549,CRC_OUT_8_27,II7547);
  nand NAND2_1463(WX2531,II7548,II7549);
  nand NAND2_1464(II7554,WX1909,CRC_OUT_8_26);
  nand NAND2_1465(II7555,WX1909,II7554);
  nand NAND2_1466(II7556,CRC_OUT_8_26,II7554);
  nand NAND2_1467(WX2532,II7555,II7556);
  nand NAND2_1468(II7561,WX1910,CRC_OUT_8_25);
  nand NAND2_1469(II7562,WX1910,II7561);
  nand NAND2_1470(II7563,CRC_OUT_8_25,II7561);
  nand NAND2_1471(WX2533,II7562,II7563);
  nand NAND2_1472(II7568,WX1911,CRC_OUT_8_24);
  nand NAND2_1473(II7569,WX1911,II7568);
  nand NAND2_1474(II7570,CRC_OUT_8_24,II7568);
  nand NAND2_1475(WX2534,II7569,II7570);
  nand NAND2_1476(II7575,WX1912,CRC_OUT_8_23);
  nand NAND2_1477(II7576,WX1912,II7575);
  nand NAND2_1478(II7577,CRC_OUT_8_23,II7575);
  nand NAND2_1479(WX2535,II7576,II7577);
  nand NAND2_1480(II7582,WX1913,CRC_OUT_8_22);
  nand NAND2_1481(II7583,WX1913,II7582);
  nand NAND2_1482(II7584,CRC_OUT_8_22,II7582);
  nand NAND2_1483(WX2536,II7583,II7584);
  nand NAND2_1484(II7589,WX1914,CRC_OUT_8_21);
  nand NAND2_1485(II7590,WX1914,II7589);
  nand NAND2_1486(II7591,CRC_OUT_8_21,II7589);
  nand NAND2_1487(WX2537,II7590,II7591);
  nand NAND2_1488(II7596,WX1915,CRC_OUT_8_20);
  nand NAND2_1489(II7597,WX1915,II7596);
  nand NAND2_1490(II7598,CRC_OUT_8_20,II7596);
  nand NAND2_1491(WX2538,II7597,II7598);
  nand NAND2_1492(II7603,WX1916,CRC_OUT_8_19);
  nand NAND2_1493(II7604,WX1916,II7603);
  nand NAND2_1494(II7605,CRC_OUT_8_19,II7603);
  nand NAND2_1495(WX2539,II7604,II7605);
  nand NAND2_1496(II7610,WX1917,CRC_OUT_8_18);
  nand NAND2_1497(II7611,WX1917,II7610);
  nand NAND2_1498(II7612,CRC_OUT_8_18,II7610);
  nand NAND2_1499(WX2540,II7611,II7612);
  nand NAND2_1500(II7617,WX1918,CRC_OUT_8_17);
  nand NAND2_1501(II7618,WX1918,II7617);
  nand NAND2_1502(II7619,CRC_OUT_8_17,II7617);
  nand NAND2_1503(WX2541,II7618,II7619);
  nand NAND2_1504(II7624,WX1919,CRC_OUT_8_16);
  nand NAND2_1505(II7625,WX1919,II7624);
  nand NAND2_1506(II7626,CRC_OUT_8_16,II7624);
  nand NAND2_1507(WX2542,II7625,II7626);
  nand NAND2_1508(II7631,WX1921,CRC_OUT_8_14);
  nand NAND2_1509(II7632,WX1921,II7631);
  nand NAND2_1510(II7633,CRC_OUT_8_14,II7631);
  nand NAND2_1511(WX2543,II7632,II7633);
  nand NAND2_1512(II7638,WX1922,CRC_OUT_8_13);
  nand NAND2_1513(II7639,WX1922,II7638);
  nand NAND2_1514(II7640,CRC_OUT_8_13,II7638);
  nand NAND2_1515(WX2544,II7639,II7640);
  nand NAND2_1516(II7645,WX1923,CRC_OUT_8_12);
  nand NAND2_1517(II7646,WX1923,II7645);
  nand NAND2_1518(II7647,CRC_OUT_8_12,II7645);
  nand NAND2_1519(WX2545,II7646,II7647);
  nand NAND2_1520(II7652,WX1924,CRC_OUT_8_11);
  nand NAND2_1521(II7653,WX1924,II7652);
  nand NAND2_1522(II7654,CRC_OUT_8_11,II7652);
  nand NAND2_1523(WX2546,II7653,II7654);
  nand NAND2_1524(II7659,WX1926,CRC_OUT_8_9);
  nand NAND2_1525(II7660,WX1926,II7659);
  nand NAND2_1526(II7661,CRC_OUT_8_9,II7659);
  nand NAND2_1527(WX2547,II7660,II7661);
  nand NAND2_1528(II7666,WX1927,CRC_OUT_8_8);
  nand NAND2_1529(II7667,WX1927,II7666);
  nand NAND2_1530(II7668,CRC_OUT_8_8,II7666);
  nand NAND2_1531(WX2548,II7667,II7668);
  nand NAND2_1532(II7673,WX1928,CRC_OUT_8_7);
  nand NAND2_1533(II7674,WX1928,II7673);
  nand NAND2_1534(II7675,CRC_OUT_8_7,II7673);
  nand NAND2_1535(WX2549,II7674,II7675);
  nand NAND2_1536(II7680,WX1929,CRC_OUT_8_6);
  nand NAND2_1537(II7681,WX1929,II7680);
  nand NAND2_1538(II7682,CRC_OUT_8_6,II7680);
  nand NAND2_1539(WX2550,II7681,II7682);
  nand NAND2_1540(II7687,WX1930,CRC_OUT_8_5);
  nand NAND2_1541(II7688,WX1930,II7687);
  nand NAND2_1542(II7689,CRC_OUT_8_5,II7687);
  nand NAND2_1543(WX2551,II7688,II7689);
  nand NAND2_1544(II7694,WX1931,CRC_OUT_8_4);
  nand NAND2_1545(II7695,WX1931,II7694);
  nand NAND2_1546(II7696,CRC_OUT_8_4,II7694);
  nand NAND2_1547(WX2552,II7695,II7696);
  nand NAND2_1548(II7701,WX1933,CRC_OUT_8_2);
  nand NAND2_1549(II7702,WX1933,II7701);
  nand NAND2_1550(II7703,CRC_OUT_8_2,II7701);
  nand NAND2_1551(WX2553,II7702,II7703);
  nand NAND2_1552(II7708,WX1934,CRC_OUT_8_1);
  nand NAND2_1553(II7709,WX1934,II7708);
  nand NAND2_1554(II7710,CRC_OUT_8_1,II7708);
  nand NAND2_1555(WX2554,II7709,II7710);
  nand NAND2_1556(II7715,WX1935,CRC_OUT_8_0);
  nand NAND2_1557(II7716,WX1935,II7715);
  nand NAND2_1558(II7717,CRC_OUT_8_0,II7715);
  nand NAND2_1559(WX2555,II7716,II7717);
  nand NAND2_1560(II9998,WX3587,WX3231);
  nand NAND2_1561(II9999,WX3587,II9998);
  nand NAND2_1562(II10000,WX3231,II9998);
  nand NAND2_1563(II9997,II9999,II10000);
  nand NAND2_1564(II10005,WX3295,II9997);
  nand NAND2_1565(II10006,WX3295,II10005);
  nand NAND2_1566(II10007,II9997,II10005);
  nand NAND2_1567(II9996,II10006,II10007);
  nand NAND2_1568(II10013,WX3359,WX3423);
  nand NAND2_1569(II10014,WX3359,II10013);
  nand NAND2_1570(II10015,WX3423,II10013);
  nand NAND2_1571(II10012,II10014,II10015);
  nand NAND2_1572(II10020,II9996,II10012);
  nand NAND2_1573(II10021,II9996,II10020);
  nand NAND2_1574(II10022,II10012,II10020);
  nand NAND2_1575(WX3486,II10021,II10022);
  nand NAND2_1576(II10029,WX3587,WX3233);
  nand NAND2_1577(II10030,WX3587,II10029);
  nand NAND2_1578(II10031,WX3233,II10029);
  nand NAND2_1579(II10028,II10030,II10031);
  nand NAND2_1580(II10036,WX3297,II10028);
  nand NAND2_1581(II10037,WX3297,II10036);
  nand NAND2_1582(II10038,II10028,II10036);
  nand NAND2_1583(II10027,II10037,II10038);
  nand NAND2_1584(II10044,WX3361,WX3425);
  nand NAND2_1585(II10045,WX3361,II10044);
  nand NAND2_1586(II10046,WX3425,II10044);
  nand NAND2_1587(II10043,II10045,II10046);
  nand NAND2_1588(II10051,II10027,II10043);
  nand NAND2_1589(II10052,II10027,II10051);
  nand NAND2_1590(II10053,II10043,II10051);
  nand NAND2_1591(WX3487,II10052,II10053);
  nand NAND2_1592(II10060,WX3587,WX3235);
  nand NAND2_1593(II10061,WX3587,II10060);
  nand NAND2_1594(II10062,WX3235,II10060);
  nand NAND2_1595(II10059,II10061,II10062);
  nand NAND2_1596(II10067,WX3299,II10059);
  nand NAND2_1597(II10068,WX3299,II10067);
  nand NAND2_1598(II10069,II10059,II10067);
  nand NAND2_1599(II10058,II10068,II10069);
  nand NAND2_1600(II10075,WX3363,WX3427);
  nand NAND2_1601(II10076,WX3363,II10075);
  nand NAND2_1602(II10077,WX3427,II10075);
  nand NAND2_1603(II10074,II10076,II10077);
  nand NAND2_1604(II10082,II10058,II10074);
  nand NAND2_1605(II10083,II10058,II10082);
  nand NAND2_1606(II10084,II10074,II10082);
  nand NAND2_1607(WX3488,II10083,II10084);
  nand NAND2_1608(II10091,WX3587,WX3237);
  nand NAND2_1609(II10092,WX3587,II10091);
  nand NAND2_1610(II10093,WX3237,II10091);
  nand NAND2_1611(II10090,II10092,II10093);
  nand NAND2_1612(II10098,WX3301,II10090);
  nand NAND2_1613(II10099,WX3301,II10098);
  nand NAND2_1614(II10100,II10090,II10098);
  nand NAND2_1615(II10089,II10099,II10100);
  nand NAND2_1616(II10106,WX3365,WX3429);
  nand NAND2_1617(II10107,WX3365,II10106);
  nand NAND2_1618(II10108,WX3429,II10106);
  nand NAND2_1619(II10105,II10107,II10108);
  nand NAND2_1620(II10113,II10089,II10105);
  nand NAND2_1621(II10114,II10089,II10113);
  nand NAND2_1622(II10115,II10105,II10113);
  nand NAND2_1623(WX3489,II10114,II10115);
  nand NAND2_1624(II10122,WX3587,WX3239);
  nand NAND2_1625(II10123,WX3587,II10122);
  nand NAND2_1626(II10124,WX3239,II10122);
  nand NAND2_1627(II10121,II10123,II10124);
  nand NAND2_1628(II10129,WX3303,II10121);
  nand NAND2_1629(II10130,WX3303,II10129);
  nand NAND2_1630(II10131,II10121,II10129);
  nand NAND2_1631(II10120,II10130,II10131);
  nand NAND2_1632(II10137,WX3367,WX3431);
  nand NAND2_1633(II10138,WX3367,II10137);
  nand NAND2_1634(II10139,WX3431,II10137);
  nand NAND2_1635(II10136,II10138,II10139);
  nand NAND2_1636(II10144,II10120,II10136);
  nand NAND2_1637(II10145,II10120,II10144);
  nand NAND2_1638(II10146,II10136,II10144);
  nand NAND2_1639(WX3490,II10145,II10146);
  nand NAND2_1640(II10153,WX3587,WX3241);
  nand NAND2_1641(II10154,WX3587,II10153);
  nand NAND2_1642(II10155,WX3241,II10153);
  nand NAND2_1643(II10152,II10154,II10155);
  nand NAND2_1644(II10160,WX3305,II10152);
  nand NAND2_1645(II10161,WX3305,II10160);
  nand NAND2_1646(II10162,II10152,II10160);
  nand NAND2_1647(II10151,II10161,II10162);
  nand NAND2_1648(II10168,WX3369,WX3433);
  nand NAND2_1649(II10169,WX3369,II10168);
  nand NAND2_1650(II10170,WX3433,II10168);
  nand NAND2_1651(II10167,II10169,II10170);
  nand NAND2_1652(II10175,II10151,II10167);
  nand NAND2_1653(II10176,II10151,II10175);
  nand NAND2_1654(II10177,II10167,II10175);
  nand NAND2_1655(WX3491,II10176,II10177);
  nand NAND2_1656(II10184,WX3587,WX3243);
  nand NAND2_1657(II10185,WX3587,II10184);
  nand NAND2_1658(II10186,WX3243,II10184);
  nand NAND2_1659(II10183,II10185,II10186);
  nand NAND2_1660(II10191,WX3307,II10183);
  nand NAND2_1661(II10192,WX3307,II10191);
  nand NAND2_1662(II10193,II10183,II10191);
  nand NAND2_1663(II10182,II10192,II10193);
  nand NAND2_1664(II10199,WX3371,WX3435);
  nand NAND2_1665(II10200,WX3371,II10199);
  nand NAND2_1666(II10201,WX3435,II10199);
  nand NAND2_1667(II10198,II10200,II10201);
  nand NAND2_1668(II10206,II10182,II10198);
  nand NAND2_1669(II10207,II10182,II10206);
  nand NAND2_1670(II10208,II10198,II10206);
  nand NAND2_1671(WX3492,II10207,II10208);
  nand NAND2_1672(II10215,WX3587,WX3245);
  nand NAND2_1673(II10216,WX3587,II10215);
  nand NAND2_1674(II10217,WX3245,II10215);
  nand NAND2_1675(II10214,II10216,II10217);
  nand NAND2_1676(II10222,WX3309,II10214);
  nand NAND2_1677(II10223,WX3309,II10222);
  nand NAND2_1678(II10224,II10214,II10222);
  nand NAND2_1679(II10213,II10223,II10224);
  nand NAND2_1680(II10230,WX3373,WX3437);
  nand NAND2_1681(II10231,WX3373,II10230);
  nand NAND2_1682(II10232,WX3437,II10230);
  nand NAND2_1683(II10229,II10231,II10232);
  nand NAND2_1684(II10237,II10213,II10229);
  nand NAND2_1685(II10238,II10213,II10237);
  nand NAND2_1686(II10239,II10229,II10237);
  nand NAND2_1687(WX3493,II10238,II10239);
  nand NAND2_1688(II10246,WX3587,WX3247);
  nand NAND2_1689(II10247,WX3587,II10246);
  nand NAND2_1690(II10248,WX3247,II10246);
  nand NAND2_1691(II10245,II10247,II10248);
  nand NAND2_1692(II10253,WX3311,II10245);
  nand NAND2_1693(II10254,WX3311,II10253);
  nand NAND2_1694(II10255,II10245,II10253);
  nand NAND2_1695(II10244,II10254,II10255);
  nand NAND2_1696(II10261,WX3375,WX3439);
  nand NAND2_1697(II10262,WX3375,II10261);
  nand NAND2_1698(II10263,WX3439,II10261);
  nand NAND2_1699(II10260,II10262,II10263);
  nand NAND2_1700(II10268,II10244,II10260);
  nand NAND2_1701(II10269,II10244,II10268);
  nand NAND2_1702(II10270,II10260,II10268);
  nand NAND2_1703(WX3494,II10269,II10270);
  nand NAND2_1704(II10277,WX3587,WX3249);
  nand NAND2_1705(II10278,WX3587,II10277);
  nand NAND2_1706(II10279,WX3249,II10277);
  nand NAND2_1707(II10276,II10278,II10279);
  nand NAND2_1708(II10284,WX3313,II10276);
  nand NAND2_1709(II10285,WX3313,II10284);
  nand NAND2_1710(II10286,II10276,II10284);
  nand NAND2_1711(II10275,II10285,II10286);
  nand NAND2_1712(II10292,WX3377,WX3441);
  nand NAND2_1713(II10293,WX3377,II10292);
  nand NAND2_1714(II10294,WX3441,II10292);
  nand NAND2_1715(II10291,II10293,II10294);
  nand NAND2_1716(II10299,II10275,II10291);
  nand NAND2_1717(II10300,II10275,II10299);
  nand NAND2_1718(II10301,II10291,II10299);
  nand NAND2_1719(WX3495,II10300,II10301);
  nand NAND2_1720(II10308,WX3587,WX3251);
  nand NAND2_1721(II10309,WX3587,II10308);
  nand NAND2_1722(II10310,WX3251,II10308);
  nand NAND2_1723(II10307,II10309,II10310);
  nand NAND2_1724(II10315,WX3315,II10307);
  nand NAND2_1725(II10316,WX3315,II10315);
  nand NAND2_1726(II10317,II10307,II10315);
  nand NAND2_1727(II10306,II10316,II10317);
  nand NAND2_1728(II10323,WX3379,WX3443);
  nand NAND2_1729(II10324,WX3379,II10323);
  nand NAND2_1730(II10325,WX3443,II10323);
  nand NAND2_1731(II10322,II10324,II10325);
  nand NAND2_1732(II10330,II10306,II10322);
  nand NAND2_1733(II10331,II10306,II10330);
  nand NAND2_1734(II10332,II10322,II10330);
  nand NAND2_1735(WX3496,II10331,II10332);
  nand NAND2_1736(II10339,WX3587,WX3253);
  nand NAND2_1737(II10340,WX3587,II10339);
  nand NAND2_1738(II10341,WX3253,II10339);
  nand NAND2_1739(II10338,II10340,II10341);
  nand NAND2_1740(II10346,WX3317,II10338);
  nand NAND2_1741(II10347,WX3317,II10346);
  nand NAND2_1742(II10348,II10338,II10346);
  nand NAND2_1743(II10337,II10347,II10348);
  nand NAND2_1744(II10354,WX3381,WX3445);
  nand NAND2_1745(II10355,WX3381,II10354);
  nand NAND2_1746(II10356,WX3445,II10354);
  nand NAND2_1747(II10353,II10355,II10356);
  nand NAND2_1748(II10361,II10337,II10353);
  nand NAND2_1749(II10362,II10337,II10361);
  nand NAND2_1750(II10363,II10353,II10361);
  nand NAND2_1751(WX3497,II10362,II10363);
  nand NAND2_1752(II10370,WX3587,WX3255);
  nand NAND2_1753(II10371,WX3587,II10370);
  nand NAND2_1754(II10372,WX3255,II10370);
  nand NAND2_1755(II10369,II10371,II10372);
  nand NAND2_1756(II10377,WX3319,II10369);
  nand NAND2_1757(II10378,WX3319,II10377);
  nand NAND2_1758(II10379,II10369,II10377);
  nand NAND2_1759(II10368,II10378,II10379);
  nand NAND2_1760(II10385,WX3383,WX3447);
  nand NAND2_1761(II10386,WX3383,II10385);
  nand NAND2_1762(II10387,WX3447,II10385);
  nand NAND2_1763(II10384,II10386,II10387);
  nand NAND2_1764(II10392,II10368,II10384);
  nand NAND2_1765(II10393,II10368,II10392);
  nand NAND2_1766(II10394,II10384,II10392);
  nand NAND2_1767(WX3498,II10393,II10394);
  nand NAND2_1768(II10401,WX3587,WX3257);
  nand NAND2_1769(II10402,WX3587,II10401);
  nand NAND2_1770(II10403,WX3257,II10401);
  nand NAND2_1771(II10400,II10402,II10403);
  nand NAND2_1772(II10408,WX3321,II10400);
  nand NAND2_1773(II10409,WX3321,II10408);
  nand NAND2_1774(II10410,II10400,II10408);
  nand NAND2_1775(II10399,II10409,II10410);
  nand NAND2_1776(II10416,WX3385,WX3449);
  nand NAND2_1777(II10417,WX3385,II10416);
  nand NAND2_1778(II10418,WX3449,II10416);
  nand NAND2_1779(II10415,II10417,II10418);
  nand NAND2_1780(II10423,II10399,II10415);
  nand NAND2_1781(II10424,II10399,II10423);
  nand NAND2_1782(II10425,II10415,II10423);
  nand NAND2_1783(WX3499,II10424,II10425);
  nand NAND2_1784(II10432,WX3587,WX3259);
  nand NAND2_1785(II10433,WX3587,II10432);
  nand NAND2_1786(II10434,WX3259,II10432);
  nand NAND2_1787(II10431,II10433,II10434);
  nand NAND2_1788(II10439,WX3323,II10431);
  nand NAND2_1789(II10440,WX3323,II10439);
  nand NAND2_1790(II10441,II10431,II10439);
  nand NAND2_1791(II10430,II10440,II10441);
  nand NAND2_1792(II10447,WX3387,WX3451);
  nand NAND2_1793(II10448,WX3387,II10447);
  nand NAND2_1794(II10449,WX3451,II10447);
  nand NAND2_1795(II10446,II10448,II10449);
  nand NAND2_1796(II10454,II10430,II10446);
  nand NAND2_1797(II10455,II10430,II10454);
  nand NAND2_1798(II10456,II10446,II10454);
  nand NAND2_1799(WX3500,II10455,II10456);
  nand NAND2_1800(II10463,WX3587,WX3261);
  nand NAND2_1801(II10464,WX3587,II10463);
  nand NAND2_1802(II10465,WX3261,II10463);
  nand NAND2_1803(II10462,II10464,II10465);
  nand NAND2_1804(II10470,WX3325,II10462);
  nand NAND2_1805(II10471,WX3325,II10470);
  nand NAND2_1806(II10472,II10462,II10470);
  nand NAND2_1807(II10461,II10471,II10472);
  nand NAND2_1808(II10478,WX3389,WX3453);
  nand NAND2_1809(II10479,WX3389,II10478);
  nand NAND2_1810(II10480,WX3453,II10478);
  nand NAND2_1811(II10477,II10479,II10480);
  nand NAND2_1812(II10485,II10461,II10477);
  nand NAND2_1813(II10486,II10461,II10485);
  nand NAND2_1814(II10487,II10477,II10485);
  nand NAND2_1815(WX3501,II10486,II10487);
  nand NAND2_1816(II10494,WX3588,WX3263);
  nand NAND2_1817(II10495,WX3588,II10494);
  nand NAND2_1818(II10496,WX3263,II10494);
  nand NAND2_1819(II10493,II10495,II10496);
  nand NAND2_1820(II10501,WX3327,II10493);
  nand NAND2_1821(II10502,WX3327,II10501);
  nand NAND2_1822(II10503,II10493,II10501);
  nand NAND2_1823(II10492,II10502,II10503);
  nand NAND2_1824(II10509,WX3391,WX3455);
  nand NAND2_1825(II10510,WX3391,II10509);
  nand NAND2_1826(II10511,WX3455,II10509);
  nand NAND2_1827(II10508,II10510,II10511);
  nand NAND2_1828(II10516,II10492,II10508);
  nand NAND2_1829(II10517,II10492,II10516);
  nand NAND2_1830(II10518,II10508,II10516);
  nand NAND2_1831(WX3502,II10517,II10518);
  nand NAND2_1832(II10525,WX3588,WX3265);
  nand NAND2_1833(II10526,WX3588,II10525);
  nand NAND2_1834(II10527,WX3265,II10525);
  nand NAND2_1835(II10524,II10526,II10527);
  nand NAND2_1836(II10532,WX3329,II10524);
  nand NAND2_1837(II10533,WX3329,II10532);
  nand NAND2_1838(II10534,II10524,II10532);
  nand NAND2_1839(II10523,II10533,II10534);
  nand NAND2_1840(II10540,WX3393,WX3457);
  nand NAND2_1841(II10541,WX3393,II10540);
  nand NAND2_1842(II10542,WX3457,II10540);
  nand NAND2_1843(II10539,II10541,II10542);
  nand NAND2_1844(II10547,II10523,II10539);
  nand NAND2_1845(II10548,II10523,II10547);
  nand NAND2_1846(II10549,II10539,II10547);
  nand NAND2_1847(WX3503,II10548,II10549);
  nand NAND2_1848(II10556,WX3588,WX3267);
  nand NAND2_1849(II10557,WX3588,II10556);
  nand NAND2_1850(II10558,WX3267,II10556);
  nand NAND2_1851(II10555,II10557,II10558);
  nand NAND2_1852(II10563,WX3331,II10555);
  nand NAND2_1853(II10564,WX3331,II10563);
  nand NAND2_1854(II10565,II10555,II10563);
  nand NAND2_1855(II10554,II10564,II10565);
  nand NAND2_1856(II10571,WX3395,WX3459);
  nand NAND2_1857(II10572,WX3395,II10571);
  nand NAND2_1858(II10573,WX3459,II10571);
  nand NAND2_1859(II10570,II10572,II10573);
  nand NAND2_1860(II10578,II10554,II10570);
  nand NAND2_1861(II10579,II10554,II10578);
  nand NAND2_1862(II10580,II10570,II10578);
  nand NAND2_1863(WX3504,II10579,II10580);
  nand NAND2_1864(II10587,WX3588,WX3269);
  nand NAND2_1865(II10588,WX3588,II10587);
  nand NAND2_1866(II10589,WX3269,II10587);
  nand NAND2_1867(II10586,II10588,II10589);
  nand NAND2_1868(II10594,WX3333,II10586);
  nand NAND2_1869(II10595,WX3333,II10594);
  nand NAND2_1870(II10596,II10586,II10594);
  nand NAND2_1871(II10585,II10595,II10596);
  nand NAND2_1872(II10602,WX3397,WX3461);
  nand NAND2_1873(II10603,WX3397,II10602);
  nand NAND2_1874(II10604,WX3461,II10602);
  nand NAND2_1875(II10601,II10603,II10604);
  nand NAND2_1876(II10609,II10585,II10601);
  nand NAND2_1877(II10610,II10585,II10609);
  nand NAND2_1878(II10611,II10601,II10609);
  nand NAND2_1879(WX3505,II10610,II10611);
  nand NAND2_1880(II10618,WX3588,WX3271);
  nand NAND2_1881(II10619,WX3588,II10618);
  nand NAND2_1882(II10620,WX3271,II10618);
  nand NAND2_1883(II10617,II10619,II10620);
  nand NAND2_1884(II10625,WX3335,II10617);
  nand NAND2_1885(II10626,WX3335,II10625);
  nand NAND2_1886(II10627,II10617,II10625);
  nand NAND2_1887(II10616,II10626,II10627);
  nand NAND2_1888(II10633,WX3399,WX3463);
  nand NAND2_1889(II10634,WX3399,II10633);
  nand NAND2_1890(II10635,WX3463,II10633);
  nand NAND2_1891(II10632,II10634,II10635);
  nand NAND2_1892(II10640,II10616,II10632);
  nand NAND2_1893(II10641,II10616,II10640);
  nand NAND2_1894(II10642,II10632,II10640);
  nand NAND2_1895(WX3506,II10641,II10642);
  nand NAND2_1896(II10649,WX3588,WX3273);
  nand NAND2_1897(II10650,WX3588,II10649);
  nand NAND2_1898(II10651,WX3273,II10649);
  nand NAND2_1899(II10648,II10650,II10651);
  nand NAND2_1900(II10656,WX3337,II10648);
  nand NAND2_1901(II10657,WX3337,II10656);
  nand NAND2_1902(II10658,II10648,II10656);
  nand NAND2_1903(II10647,II10657,II10658);
  nand NAND2_1904(II10664,WX3401,WX3465);
  nand NAND2_1905(II10665,WX3401,II10664);
  nand NAND2_1906(II10666,WX3465,II10664);
  nand NAND2_1907(II10663,II10665,II10666);
  nand NAND2_1908(II10671,II10647,II10663);
  nand NAND2_1909(II10672,II10647,II10671);
  nand NAND2_1910(II10673,II10663,II10671);
  nand NAND2_1911(WX3507,II10672,II10673);
  nand NAND2_1912(II10680,WX3588,WX3275);
  nand NAND2_1913(II10681,WX3588,II10680);
  nand NAND2_1914(II10682,WX3275,II10680);
  nand NAND2_1915(II10679,II10681,II10682);
  nand NAND2_1916(II10687,WX3339,II10679);
  nand NAND2_1917(II10688,WX3339,II10687);
  nand NAND2_1918(II10689,II10679,II10687);
  nand NAND2_1919(II10678,II10688,II10689);
  nand NAND2_1920(II10695,WX3403,WX3467);
  nand NAND2_1921(II10696,WX3403,II10695);
  nand NAND2_1922(II10697,WX3467,II10695);
  nand NAND2_1923(II10694,II10696,II10697);
  nand NAND2_1924(II10702,II10678,II10694);
  nand NAND2_1925(II10703,II10678,II10702);
  nand NAND2_1926(II10704,II10694,II10702);
  nand NAND2_1927(WX3508,II10703,II10704);
  nand NAND2_1928(II10711,WX3588,WX3277);
  nand NAND2_1929(II10712,WX3588,II10711);
  nand NAND2_1930(II10713,WX3277,II10711);
  nand NAND2_1931(II10710,II10712,II10713);
  nand NAND2_1932(II10718,WX3341,II10710);
  nand NAND2_1933(II10719,WX3341,II10718);
  nand NAND2_1934(II10720,II10710,II10718);
  nand NAND2_1935(II10709,II10719,II10720);
  nand NAND2_1936(II10726,WX3405,WX3469);
  nand NAND2_1937(II10727,WX3405,II10726);
  nand NAND2_1938(II10728,WX3469,II10726);
  nand NAND2_1939(II10725,II10727,II10728);
  nand NAND2_1940(II10733,II10709,II10725);
  nand NAND2_1941(II10734,II10709,II10733);
  nand NAND2_1942(II10735,II10725,II10733);
  nand NAND2_1943(WX3509,II10734,II10735);
  nand NAND2_1944(II10742,WX3588,WX3279);
  nand NAND2_1945(II10743,WX3588,II10742);
  nand NAND2_1946(II10744,WX3279,II10742);
  nand NAND2_1947(II10741,II10743,II10744);
  nand NAND2_1948(II10749,WX3343,II10741);
  nand NAND2_1949(II10750,WX3343,II10749);
  nand NAND2_1950(II10751,II10741,II10749);
  nand NAND2_1951(II10740,II10750,II10751);
  nand NAND2_1952(II10757,WX3407,WX3471);
  nand NAND2_1953(II10758,WX3407,II10757);
  nand NAND2_1954(II10759,WX3471,II10757);
  nand NAND2_1955(II10756,II10758,II10759);
  nand NAND2_1956(II10764,II10740,II10756);
  nand NAND2_1957(II10765,II10740,II10764);
  nand NAND2_1958(II10766,II10756,II10764);
  nand NAND2_1959(WX3510,II10765,II10766);
  nand NAND2_1960(II10773,WX3588,WX3281);
  nand NAND2_1961(II10774,WX3588,II10773);
  nand NAND2_1962(II10775,WX3281,II10773);
  nand NAND2_1963(II10772,II10774,II10775);
  nand NAND2_1964(II10780,WX3345,II10772);
  nand NAND2_1965(II10781,WX3345,II10780);
  nand NAND2_1966(II10782,II10772,II10780);
  nand NAND2_1967(II10771,II10781,II10782);
  nand NAND2_1968(II10788,WX3409,WX3473);
  nand NAND2_1969(II10789,WX3409,II10788);
  nand NAND2_1970(II10790,WX3473,II10788);
  nand NAND2_1971(II10787,II10789,II10790);
  nand NAND2_1972(II10795,II10771,II10787);
  nand NAND2_1973(II10796,II10771,II10795);
  nand NAND2_1974(II10797,II10787,II10795);
  nand NAND2_1975(WX3511,II10796,II10797);
  nand NAND2_1976(II10804,WX3588,WX3283);
  nand NAND2_1977(II10805,WX3588,II10804);
  nand NAND2_1978(II10806,WX3283,II10804);
  nand NAND2_1979(II10803,II10805,II10806);
  nand NAND2_1980(II10811,WX3347,II10803);
  nand NAND2_1981(II10812,WX3347,II10811);
  nand NAND2_1982(II10813,II10803,II10811);
  nand NAND2_1983(II10802,II10812,II10813);
  nand NAND2_1984(II10819,WX3411,WX3475);
  nand NAND2_1985(II10820,WX3411,II10819);
  nand NAND2_1986(II10821,WX3475,II10819);
  nand NAND2_1987(II10818,II10820,II10821);
  nand NAND2_1988(II10826,II10802,II10818);
  nand NAND2_1989(II10827,II10802,II10826);
  nand NAND2_1990(II10828,II10818,II10826);
  nand NAND2_1991(WX3512,II10827,II10828);
  nand NAND2_1992(II10835,WX3588,WX3285);
  nand NAND2_1993(II10836,WX3588,II10835);
  nand NAND2_1994(II10837,WX3285,II10835);
  nand NAND2_1995(II10834,II10836,II10837);
  nand NAND2_1996(II10842,WX3349,II10834);
  nand NAND2_1997(II10843,WX3349,II10842);
  nand NAND2_1998(II10844,II10834,II10842);
  nand NAND2_1999(II10833,II10843,II10844);
  nand NAND2_2000(II10850,WX3413,WX3477);
  nand NAND2_2001(II10851,WX3413,II10850);
  nand NAND2_2002(II10852,WX3477,II10850);
  nand NAND2_2003(II10849,II10851,II10852);
  nand NAND2_2004(II10857,II10833,II10849);
  nand NAND2_2005(II10858,II10833,II10857);
  nand NAND2_2006(II10859,II10849,II10857);
  nand NAND2_2007(WX3513,II10858,II10859);
  nand NAND2_2008(II10866,WX3588,WX3287);
  nand NAND2_2009(II10867,WX3588,II10866);
  nand NAND2_2010(II10868,WX3287,II10866);
  nand NAND2_2011(II10865,II10867,II10868);
  nand NAND2_2012(II10873,WX3351,II10865);
  nand NAND2_2013(II10874,WX3351,II10873);
  nand NAND2_2014(II10875,II10865,II10873);
  nand NAND2_2015(II10864,II10874,II10875);
  nand NAND2_2016(II10881,WX3415,WX3479);
  nand NAND2_2017(II10882,WX3415,II10881);
  nand NAND2_2018(II10883,WX3479,II10881);
  nand NAND2_2019(II10880,II10882,II10883);
  nand NAND2_2020(II10888,II10864,II10880);
  nand NAND2_2021(II10889,II10864,II10888);
  nand NAND2_2022(II10890,II10880,II10888);
  nand NAND2_2023(WX3514,II10889,II10890);
  nand NAND2_2024(II10897,WX3588,WX3289);
  nand NAND2_2025(II10898,WX3588,II10897);
  nand NAND2_2026(II10899,WX3289,II10897);
  nand NAND2_2027(II10896,II10898,II10899);
  nand NAND2_2028(II10904,WX3353,II10896);
  nand NAND2_2029(II10905,WX3353,II10904);
  nand NAND2_2030(II10906,II10896,II10904);
  nand NAND2_2031(II10895,II10905,II10906);
  nand NAND2_2032(II10912,WX3417,WX3481);
  nand NAND2_2033(II10913,WX3417,II10912);
  nand NAND2_2034(II10914,WX3481,II10912);
  nand NAND2_2035(II10911,II10913,II10914);
  nand NAND2_2036(II10919,II10895,II10911);
  nand NAND2_2037(II10920,II10895,II10919);
  nand NAND2_2038(II10921,II10911,II10919);
  nand NAND2_2039(WX3515,II10920,II10921);
  nand NAND2_2040(II10928,WX3588,WX3291);
  nand NAND2_2041(II10929,WX3588,II10928);
  nand NAND2_2042(II10930,WX3291,II10928);
  nand NAND2_2043(II10927,II10929,II10930);
  nand NAND2_2044(II10935,WX3355,II10927);
  nand NAND2_2045(II10936,WX3355,II10935);
  nand NAND2_2046(II10937,II10927,II10935);
  nand NAND2_2047(II10926,II10936,II10937);
  nand NAND2_2048(II10943,WX3419,WX3483);
  nand NAND2_2049(II10944,WX3419,II10943);
  nand NAND2_2050(II10945,WX3483,II10943);
  nand NAND2_2051(II10942,II10944,II10945);
  nand NAND2_2052(II10950,II10926,II10942);
  nand NAND2_2053(II10951,II10926,II10950);
  nand NAND2_2054(II10952,II10942,II10950);
  nand NAND2_2055(WX3516,II10951,II10952);
  nand NAND2_2056(II10959,WX3588,WX3293);
  nand NAND2_2057(II10960,WX3588,II10959);
  nand NAND2_2058(II10961,WX3293,II10959);
  nand NAND2_2059(II10958,II10960,II10961);
  nand NAND2_2060(II10966,WX3357,II10958);
  nand NAND2_2061(II10967,WX3357,II10966);
  nand NAND2_2062(II10968,II10958,II10966);
  nand NAND2_2063(II10957,II10967,II10968);
  nand NAND2_2064(II10974,WX3421,WX3485);
  nand NAND2_2065(II10975,WX3421,II10974);
  nand NAND2_2066(II10976,WX3485,II10974);
  nand NAND2_2067(II10973,II10975,II10976);
  nand NAND2_2068(II10981,II10957,II10973);
  nand NAND2_2069(II10982,II10957,II10981);
  nand NAND2_2070(II10983,II10973,II10981);
  nand NAND2_2071(WX3517,II10982,II10983);
  nand NAND2_2072(II11062,WX3166,WX3071);
  nand NAND2_2073(II11063,WX3166,II11062);
  nand NAND2_2074(II11064,WX3071,II11062);
  nand NAND2_2075(WX3592,II11063,II11064);
  nand NAND2_2076(II11075,WX3167,WX3073);
  nand NAND2_2077(II11076,WX3167,II11075);
  nand NAND2_2078(II11077,WX3073,II11075);
  nand NAND2_2079(WX3599,II11076,II11077);
  nand NAND2_2080(II11088,WX3168,WX3075);
  nand NAND2_2081(II11089,WX3168,II11088);
  nand NAND2_2082(II11090,WX3075,II11088);
  nand NAND2_2083(WX3606,II11089,II11090);
  nand NAND2_2084(II11101,WX3169,WX3077);
  nand NAND2_2085(II11102,WX3169,II11101);
  nand NAND2_2086(II11103,WX3077,II11101);
  nand NAND2_2087(WX3613,II11102,II11103);
  nand NAND2_2088(II11114,WX3170,WX3079);
  nand NAND2_2089(II11115,WX3170,II11114);
  nand NAND2_2090(II11116,WX3079,II11114);
  nand NAND2_2091(WX3620,II11115,II11116);
  nand NAND2_2092(II11127,WX3171,WX3081);
  nand NAND2_2093(II11128,WX3171,II11127);
  nand NAND2_2094(II11129,WX3081,II11127);
  nand NAND2_2095(WX3627,II11128,II11129);
  nand NAND2_2096(II11140,WX3172,WX3083);
  nand NAND2_2097(II11141,WX3172,II11140);
  nand NAND2_2098(II11142,WX3083,II11140);
  nand NAND2_2099(WX3634,II11141,II11142);
  nand NAND2_2100(II11153,WX3173,WX3085);
  nand NAND2_2101(II11154,WX3173,II11153);
  nand NAND2_2102(II11155,WX3085,II11153);
  nand NAND2_2103(WX3641,II11154,II11155);
  nand NAND2_2104(II11166,WX3174,WX3087);
  nand NAND2_2105(II11167,WX3174,II11166);
  nand NAND2_2106(II11168,WX3087,II11166);
  nand NAND2_2107(WX3648,II11167,II11168);
  nand NAND2_2108(II11179,WX3175,WX3089);
  nand NAND2_2109(II11180,WX3175,II11179);
  nand NAND2_2110(II11181,WX3089,II11179);
  nand NAND2_2111(WX3655,II11180,II11181);
  nand NAND2_2112(II11192,WX3176,WX3091);
  nand NAND2_2113(II11193,WX3176,II11192);
  nand NAND2_2114(II11194,WX3091,II11192);
  nand NAND2_2115(WX3662,II11193,II11194);
  nand NAND2_2116(II11205,WX3177,WX3093);
  nand NAND2_2117(II11206,WX3177,II11205);
  nand NAND2_2118(II11207,WX3093,II11205);
  nand NAND2_2119(WX3669,II11206,II11207);
  nand NAND2_2120(II11218,WX3178,WX3095);
  nand NAND2_2121(II11219,WX3178,II11218);
  nand NAND2_2122(II11220,WX3095,II11218);
  nand NAND2_2123(WX3676,II11219,II11220);
  nand NAND2_2124(II11231,WX3179,WX3097);
  nand NAND2_2125(II11232,WX3179,II11231);
  nand NAND2_2126(II11233,WX3097,II11231);
  nand NAND2_2127(WX3683,II11232,II11233);
  nand NAND2_2128(II11244,WX3180,WX3099);
  nand NAND2_2129(II11245,WX3180,II11244);
  nand NAND2_2130(II11246,WX3099,II11244);
  nand NAND2_2131(WX3690,II11245,II11246);
  nand NAND2_2132(II11257,WX3181,WX3101);
  nand NAND2_2133(II11258,WX3181,II11257);
  nand NAND2_2134(II11259,WX3101,II11257);
  nand NAND2_2135(WX3697,II11258,II11259);
  nand NAND2_2136(II11270,WX3182,WX3103);
  nand NAND2_2137(II11271,WX3182,II11270);
  nand NAND2_2138(II11272,WX3103,II11270);
  nand NAND2_2139(WX3704,II11271,II11272);
  nand NAND2_2140(II11283,WX3183,WX3105);
  nand NAND2_2141(II11284,WX3183,II11283);
  nand NAND2_2142(II11285,WX3105,II11283);
  nand NAND2_2143(WX3711,II11284,II11285);
  nand NAND2_2144(II11296,WX3184,WX3107);
  nand NAND2_2145(II11297,WX3184,II11296);
  nand NAND2_2146(II11298,WX3107,II11296);
  nand NAND2_2147(WX3718,II11297,II11298);
  nand NAND2_2148(II11309,WX3185,WX3109);
  nand NAND2_2149(II11310,WX3185,II11309);
  nand NAND2_2150(II11311,WX3109,II11309);
  nand NAND2_2151(WX3725,II11310,II11311);
  nand NAND2_2152(II11322,WX3186,WX3111);
  nand NAND2_2153(II11323,WX3186,II11322);
  nand NAND2_2154(II11324,WX3111,II11322);
  nand NAND2_2155(WX3732,II11323,II11324);
  nand NAND2_2156(II11335,WX3187,WX3113);
  nand NAND2_2157(II11336,WX3187,II11335);
  nand NAND2_2158(II11337,WX3113,II11335);
  nand NAND2_2159(WX3739,II11336,II11337);
  nand NAND2_2160(II11348,WX3188,WX3115);
  nand NAND2_2161(II11349,WX3188,II11348);
  nand NAND2_2162(II11350,WX3115,II11348);
  nand NAND2_2163(WX3746,II11349,II11350);
  nand NAND2_2164(II11361,WX3189,WX3117);
  nand NAND2_2165(II11362,WX3189,II11361);
  nand NAND2_2166(II11363,WX3117,II11361);
  nand NAND2_2167(WX3753,II11362,II11363);
  nand NAND2_2168(II11374,WX3190,WX3119);
  nand NAND2_2169(II11375,WX3190,II11374);
  nand NAND2_2170(II11376,WX3119,II11374);
  nand NAND2_2171(WX3760,II11375,II11376);
  nand NAND2_2172(II11387,WX3191,WX3121);
  nand NAND2_2173(II11388,WX3191,II11387);
  nand NAND2_2174(II11389,WX3121,II11387);
  nand NAND2_2175(WX3767,II11388,II11389);
  nand NAND2_2176(II11400,WX3192,WX3123);
  nand NAND2_2177(II11401,WX3192,II11400);
  nand NAND2_2178(II11402,WX3123,II11400);
  nand NAND2_2179(WX3774,II11401,II11402);
  nand NAND2_2180(II11413,WX3193,WX3125);
  nand NAND2_2181(II11414,WX3193,II11413);
  nand NAND2_2182(II11415,WX3125,II11413);
  nand NAND2_2183(WX3781,II11414,II11415);
  nand NAND2_2184(II11426,WX3194,WX3127);
  nand NAND2_2185(II11427,WX3194,II11426);
  nand NAND2_2186(II11428,WX3127,II11426);
  nand NAND2_2187(WX3788,II11427,II11428);
  nand NAND2_2188(II11439,WX3195,WX3129);
  nand NAND2_2189(II11440,WX3195,II11439);
  nand NAND2_2190(II11441,WX3129,II11439);
  nand NAND2_2191(WX3795,II11440,II11441);
  nand NAND2_2192(II11452,WX3196,WX3131);
  nand NAND2_2193(II11453,WX3196,II11452);
  nand NAND2_2194(II11454,WX3131,II11452);
  nand NAND2_2195(WX3802,II11453,II11454);
  nand NAND2_2196(II11465,WX3197,WX3133);
  nand NAND2_2197(II11466,WX3197,II11465);
  nand NAND2_2198(II11467,WX3133,II11465);
  nand NAND2_2199(WX3809,II11466,II11467);
  nand NAND2_2200(II11480,WX3213,CRC_OUT_7_31);
  nand NAND2_2201(II11481,WX3213,II11480);
  nand NAND2_2202(II11482,CRC_OUT_7_31,II11480);
  nand NAND2_2203(II11479,II11481,II11482);
  nand NAND2_2204(II11487,CRC_OUT_7_15,II11479);
  nand NAND2_2205(II11488,CRC_OUT_7_15,II11487);
  nand NAND2_2206(II11489,II11479,II11487);
  nand NAND2_2207(WX3817,II11488,II11489);
  nand NAND2_2208(II11495,WX3218,CRC_OUT_7_31);
  nand NAND2_2209(II11496,WX3218,II11495);
  nand NAND2_2210(II11497,CRC_OUT_7_31,II11495);
  nand NAND2_2211(II11494,II11496,II11497);
  nand NAND2_2212(II11502,CRC_OUT_7_10,II11494);
  nand NAND2_2213(II11503,CRC_OUT_7_10,II11502);
  nand NAND2_2214(II11504,II11494,II11502);
  nand NAND2_2215(WX3818,II11503,II11504);
  nand NAND2_2216(II11510,WX3225,CRC_OUT_7_31);
  nand NAND2_2217(II11511,WX3225,II11510);
  nand NAND2_2218(II11512,CRC_OUT_7_31,II11510);
  nand NAND2_2219(II11509,II11511,II11512);
  nand NAND2_2220(II11517,CRC_OUT_7_3,II11509);
  nand NAND2_2221(II11518,CRC_OUT_7_3,II11517);
  nand NAND2_2222(II11519,II11509,II11517);
  nand NAND2_2223(WX3819,II11518,II11519);
  nand NAND2_2224(II11524,WX3229,CRC_OUT_7_31);
  nand NAND2_2225(II11525,WX3229,II11524);
  nand NAND2_2226(II11526,CRC_OUT_7_31,II11524);
  nand NAND2_2227(WX3820,II11525,II11526);
  nand NAND2_2228(II11531,WX3198,CRC_OUT_7_30);
  nand NAND2_2229(II11532,WX3198,II11531);
  nand NAND2_2230(II11533,CRC_OUT_7_30,II11531);
  nand NAND2_2231(WX3821,II11532,II11533);
  nand NAND2_2232(II11538,WX3199,CRC_OUT_7_29);
  nand NAND2_2233(II11539,WX3199,II11538);
  nand NAND2_2234(II11540,CRC_OUT_7_29,II11538);
  nand NAND2_2235(WX3822,II11539,II11540);
  nand NAND2_2236(II11545,WX3200,CRC_OUT_7_28);
  nand NAND2_2237(II11546,WX3200,II11545);
  nand NAND2_2238(II11547,CRC_OUT_7_28,II11545);
  nand NAND2_2239(WX3823,II11546,II11547);
  nand NAND2_2240(II11552,WX3201,CRC_OUT_7_27);
  nand NAND2_2241(II11553,WX3201,II11552);
  nand NAND2_2242(II11554,CRC_OUT_7_27,II11552);
  nand NAND2_2243(WX3824,II11553,II11554);
  nand NAND2_2244(II11559,WX3202,CRC_OUT_7_26);
  nand NAND2_2245(II11560,WX3202,II11559);
  nand NAND2_2246(II11561,CRC_OUT_7_26,II11559);
  nand NAND2_2247(WX3825,II11560,II11561);
  nand NAND2_2248(II11566,WX3203,CRC_OUT_7_25);
  nand NAND2_2249(II11567,WX3203,II11566);
  nand NAND2_2250(II11568,CRC_OUT_7_25,II11566);
  nand NAND2_2251(WX3826,II11567,II11568);
  nand NAND2_2252(II11573,WX3204,CRC_OUT_7_24);
  nand NAND2_2253(II11574,WX3204,II11573);
  nand NAND2_2254(II11575,CRC_OUT_7_24,II11573);
  nand NAND2_2255(WX3827,II11574,II11575);
  nand NAND2_2256(II11580,WX3205,CRC_OUT_7_23);
  nand NAND2_2257(II11581,WX3205,II11580);
  nand NAND2_2258(II11582,CRC_OUT_7_23,II11580);
  nand NAND2_2259(WX3828,II11581,II11582);
  nand NAND2_2260(II11587,WX3206,CRC_OUT_7_22);
  nand NAND2_2261(II11588,WX3206,II11587);
  nand NAND2_2262(II11589,CRC_OUT_7_22,II11587);
  nand NAND2_2263(WX3829,II11588,II11589);
  nand NAND2_2264(II11594,WX3207,CRC_OUT_7_21);
  nand NAND2_2265(II11595,WX3207,II11594);
  nand NAND2_2266(II11596,CRC_OUT_7_21,II11594);
  nand NAND2_2267(WX3830,II11595,II11596);
  nand NAND2_2268(II11601,WX3208,CRC_OUT_7_20);
  nand NAND2_2269(II11602,WX3208,II11601);
  nand NAND2_2270(II11603,CRC_OUT_7_20,II11601);
  nand NAND2_2271(WX3831,II11602,II11603);
  nand NAND2_2272(II11608,WX3209,CRC_OUT_7_19);
  nand NAND2_2273(II11609,WX3209,II11608);
  nand NAND2_2274(II11610,CRC_OUT_7_19,II11608);
  nand NAND2_2275(WX3832,II11609,II11610);
  nand NAND2_2276(II11615,WX3210,CRC_OUT_7_18);
  nand NAND2_2277(II11616,WX3210,II11615);
  nand NAND2_2278(II11617,CRC_OUT_7_18,II11615);
  nand NAND2_2279(WX3833,II11616,II11617);
  nand NAND2_2280(II11622,WX3211,CRC_OUT_7_17);
  nand NAND2_2281(II11623,WX3211,II11622);
  nand NAND2_2282(II11624,CRC_OUT_7_17,II11622);
  nand NAND2_2283(WX3834,II11623,II11624);
  nand NAND2_2284(II11629,WX3212,CRC_OUT_7_16);
  nand NAND2_2285(II11630,WX3212,II11629);
  nand NAND2_2286(II11631,CRC_OUT_7_16,II11629);
  nand NAND2_2287(WX3835,II11630,II11631);
  nand NAND2_2288(II11636,WX3214,CRC_OUT_7_14);
  nand NAND2_2289(II11637,WX3214,II11636);
  nand NAND2_2290(II11638,CRC_OUT_7_14,II11636);
  nand NAND2_2291(WX3836,II11637,II11638);
  nand NAND2_2292(II11643,WX3215,CRC_OUT_7_13);
  nand NAND2_2293(II11644,WX3215,II11643);
  nand NAND2_2294(II11645,CRC_OUT_7_13,II11643);
  nand NAND2_2295(WX3837,II11644,II11645);
  nand NAND2_2296(II11650,WX3216,CRC_OUT_7_12);
  nand NAND2_2297(II11651,WX3216,II11650);
  nand NAND2_2298(II11652,CRC_OUT_7_12,II11650);
  nand NAND2_2299(WX3838,II11651,II11652);
  nand NAND2_2300(II11657,WX3217,CRC_OUT_7_11);
  nand NAND2_2301(II11658,WX3217,II11657);
  nand NAND2_2302(II11659,CRC_OUT_7_11,II11657);
  nand NAND2_2303(WX3839,II11658,II11659);
  nand NAND2_2304(II11664,WX3219,CRC_OUT_7_9);
  nand NAND2_2305(II11665,WX3219,II11664);
  nand NAND2_2306(II11666,CRC_OUT_7_9,II11664);
  nand NAND2_2307(WX3840,II11665,II11666);
  nand NAND2_2308(II11671,WX3220,CRC_OUT_7_8);
  nand NAND2_2309(II11672,WX3220,II11671);
  nand NAND2_2310(II11673,CRC_OUT_7_8,II11671);
  nand NAND2_2311(WX3841,II11672,II11673);
  nand NAND2_2312(II11678,WX3221,CRC_OUT_7_7);
  nand NAND2_2313(II11679,WX3221,II11678);
  nand NAND2_2314(II11680,CRC_OUT_7_7,II11678);
  nand NAND2_2315(WX3842,II11679,II11680);
  nand NAND2_2316(II11685,WX3222,CRC_OUT_7_6);
  nand NAND2_2317(II11686,WX3222,II11685);
  nand NAND2_2318(II11687,CRC_OUT_7_6,II11685);
  nand NAND2_2319(WX3843,II11686,II11687);
  nand NAND2_2320(II11692,WX3223,CRC_OUT_7_5);
  nand NAND2_2321(II11693,WX3223,II11692);
  nand NAND2_2322(II11694,CRC_OUT_7_5,II11692);
  nand NAND2_2323(WX3844,II11693,II11694);
  nand NAND2_2324(II11699,WX3224,CRC_OUT_7_4);
  nand NAND2_2325(II11700,WX3224,II11699);
  nand NAND2_2326(II11701,CRC_OUT_7_4,II11699);
  nand NAND2_2327(WX3845,II11700,II11701);
  nand NAND2_2328(II11706,WX3226,CRC_OUT_7_2);
  nand NAND2_2329(II11707,WX3226,II11706);
  nand NAND2_2330(II11708,CRC_OUT_7_2,II11706);
  nand NAND2_2331(WX3846,II11707,II11708);
  nand NAND2_2332(II11713,WX3227,CRC_OUT_7_1);
  nand NAND2_2333(II11714,WX3227,II11713);
  nand NAND2_2334(II11715,CRC_OUT_7_1,II11713);
  nand NAND2_2335(WX3847,II11714,II11715);
  nand NAND2_2336(II11720,WX3228,CRC_OUT_7_0);
  nand NAND2_2337(II11721,WX3228,II11720);
  nand NAND2_2338(II11722,CRC_OUT_7_0,II11720);
  nand NAND2_2339(WX3848,II11721,II11722);
  nand NAND2_2340(II14003,WX4880,WX4524);
  nand NAND2_2341(II14004,WX4880,II14003);
  nand NAND2_2342(II14005,WX4524,II14003);
  nand NAND2_2343(II14002,II14004,II14005);
  nand NAND2_2344(II14010,WX4588,II14002);
  nand NAND2_2345(II14011,WX4588,II14010);
  nand NAND2_2346(II14012,II14002,II14010);
  nand NAND2_2347(II14001,II14011,II14012);
  nand NAND2_2348(II14018,WX4652,WX4716);
  nand NAND2_2349(II14019,WX4652,II14018);
  nand NAND2_2350(II14020,WX4716,II14018);
  nand NAND2_2351(II14017,II14019,II14020);
  nand NAND2_2352(II14025,II14001,II14017);
  nand NAND2_2353(II14026,II14001,II14025);
  nand NAND2_2354(II14027,II14017,II14025);
  nand NAND2_2355(WX4779,II14026,II14027);
  nand NAND2_2356(II14034,WX4880,WX4526);
  nand NAND2_2357(II14035,WX4880,II14034);
  nand NAND2_2358(II14036,WX4526,II14034);
  nand NAND2_2359(II14033,II14035,II14036);
  nand NAND2_2360(II14041,WX4590,II14033);
  nand NAND2_2361(II14042,WX4590,II14041);
  nand NAND2_2362(II14043,II14033,II14041);
  nand NAND2_2363(II14032,II14042,II14043);
  nand NAND2_2364(II14049,WX4654,WX4718);
  nand NAND2_2365(II14050,WX4654,II14049);
  nand NAND2_2366(II14051,WX4718,II14049);
  nand NAND2_2367(II14048,II14050,II14051);
  nand NAND2_2368(II14056,II14032,II14048);
  nand NAND2_2369(II14057,II14032,II14056);
  nand NAND2_2370(II14058,II14048,II14056);
  nand NAND2_2371(WX4780,II14057,II14058);
  nand NAND2_2372(II14065,WX4880,WX4528);
  nand NAND2_2373(II14066,WX4880,II14065);
  nand NAND2_2374(II14067,WX4528,II14065);
  nand NAND2_2375(II14064,II14066,II14067);
  nand NAND2_2376(II14072,WX4592,II14064);
  nand NAND2_2377(II14073,WX4592,II14072);
  nand NAND2_2378(II14074,II14064,II14072);
  nand NAND2_2379(II14063,II14073,II14074);
  nand NAND2_2380(II14080,WX4656,WX4720);
  nand NAND2_2381(II14081,WX4656,II14080);
  nand NAND2_2382(II14082,WX4720,II14080);
  nand NAND2_2383(II14079,II14081,II14082);
  nand NAND2_2384(II14087,II14063,II14079);
  nand NAND2_2385(II14088,II14063,II14087);
  nand NAND2_2386(II14089,II14079,II14087);
  nand NAND2_2387(WX4781,II14088,II14089);
  nand NAND2_2388(II14096,WX4880,WX4530);
  nand NAND2_2389(II14097,WX4880,II14096);
  nand NAND2_2390(II14098,WX4530,II14096);
  nand NAND2_2391(II14095,II14097,II14098);
  nand NAND2_2392(II14103,WX4594,II14095);
  nand NAND2_2393(II14104,WX4594,II14103);
  nand NAND2_2394(II14105,II14095,II14103);
  nand NAND2_2395(II14094,II14104,II14105);
  nand NAND2_2396(II14111,WX4658,WX4722);
  nand NAND2_2397(II14112,WX4658,II14111);
  nand NAND2_2398(II14113,WX4722,II14111);
  nand NAND2_2399(II14110,II14112,II14113);
  nand NAND2_2400(II14118,II14094,II14110);
  nand NAND2_2401(II14119,II14094,II14118);
  nand NAND2_2402(II14120,II14110,II14118);
  nand NAND2_2403(WX4782,II14119,II14120);
  nand NAND2_2404(II14127,WX4880,WX4532);
  nand NAND2_2405(II14128,WX4880,II14127);
  nand NAND2_2406(II14129,WX4532,II14127);
  nand NAND2_2407(II14126,II14128,II14129);
  nand NAND2_2408(II14134,WX4596,II14126);
  nand NAND2_2409(II14135,WX4596,II14134);
  nand NAND2_2410(II14136,II14126,II14134);
  nand NAND2_2411(II14125,II14135,II14136);
  nand NAND2_2412(II14142,WX4660,WX4724);
  nand NAND2_2413(II14143,WX4660,II14142);
  nand NAND2_2414(II14144,WX4724,II14142);
  nand NAND2_2415(II14141,II14143,II14144);
  nand NAND2_2416(II14149,II14125,II14141);
  nand NAND2_2417(II14150,II14125,II14149);
  nand NAND2_2418(II14151,II14141,II14149);
  nand NAND2_2419(WX4783,II14150,II14151);
  nand NAND2_2420(II14158,WX4880,WX4534);
  nand NAND2_2421(II14159,WX4880,II14158);
  nand NAND2_2422(II14160,WX4534,II14158);
  nand NAND2_2423(II14157,II14159,II14160);
  nand NAND2_2424(II14165,WX4598,II14157);
  nand NAND2_2425(II14166,WX4598,II14165);
  nand NAND2_2426(II14167,II14157,II14165);
  nand NAND2_2427(II14156,II14166,II14167);
  nand NAND2_2428(II14173,WX4662,WX4726);
  nand NAND2_2429(II14174,WX4662,II14173);
  nand NAND2_2430(II14175,WX4726,II14173);
  nand NAND2_2431(II14172,II14174,II14175);
  nand NAND2_2432(II14180,II14156,II14172);
  nand NAND2_2433(II14181,II14156,II14180);
  nand NAND2_2434(II14182,II14172,II14180);
  nand NAND2_2435(WX4784,II14181,II14182);
  nand NAND2_2436(II14189,WX4880,WX4536);
  nand NAND2_2437(II14190,WX4880,II14189);
  nand NAND2_2438(II14191,WX4536,II14189);
  nand NAND2_2439(II14188,II14190,II14191);
  nand NAND2_2440(II14196,WX4600,II14188);
  nand NAND2_2441(II14197,WX4600,II14196);
  nand NAND2_2442(II14198,II14188,II14196);
  nand NAND2_2443(II14187,II14197,II14198);
  nand NAND2_2444(II14204,WX4664,WX4728);
  nand NAND2_2445(II14205,WX4664,II14204);
  nand NAND2_2446(II14206,WX4728,II14204);
  nand NAND2_2447(II14203,II14205,II14206);
  nand NAND2_2448(II14211,II14187,II14203);
  nand NAND2_2449(II14212,II14187,II14211);
  nand NAND2_2450(II14213,II14203,II14211);
  nand NAND2_2451(WX4785,II14212,II14213);
  nand NAND2_2452(II14220,WX4880,WX4538);
  nand NAND2_2453(II14221,WX4880,II14220);
  nand NAND2_2454(II14222,WX4538,II14220);
  nand NAND2_2455(II14219,II14221,II14222);
  nand NAND2_2456(II14227,WX4602,II14219);
  nand NAND2_2457(II14228,WX4602,II14227);
  nand NAND2_2458(II14229,II14219,II14227);
  nand NAND2_2459(II14218,II14228,II14229);
  nand NAND2_2460(II14235,WX4666,WX4730);
  nand NAND2_2461(II14236,WX4666,II14235);
  nand NAND2_2462(II14237,WX4730,II14235);
  nand NAND2_2463(II14234,II14236,II14237);
  nand NAND2_2464(II14242,II14218,II14234);
  nand NAND2_2465(II14243,II14218,II14242);
  nand NAND2_2466(II14244,II14234,II14242);
  nand NAND2_2467(WX4786,II14243,II14244);
  nand NAND2_2468(II14251,WX4880,WX4540);
  nand NAND2_2469(II14252,WX4880,II14251);
  nand NAND2_2470(II14253,WX4540,II14251);
  nand NAND2_2471(II14250,II14252,II14253);
  nand NAND2_2472(II14258,WX4604,II14250);
  nand NAND2_2473(II14259,WX4604,II14258);
  nand NAND2_2474(II14260,II14250,II14258);
  nand NAND2_2475(II14249,II14259,II14260);
  nand NAND2_2476(II14266,WX4668,WX4732);
  nand NAND2_2477(II14267,WX4668,II14266);
  nand NAND2_2478(II14268,WX4732,II14266);
  nand NAND2_2479(II14265,II14267,II14268);
  nand NAND2_2480(II14273,II14249,II14265);
  nand NAND2_2481(II14274,II14249,II14273);
  nand NAND2_2482(II14275,II14265,II14273);
  nand NAND2_2483(WX4787,II14274,II14275);
  nand NAND2_2484(II14282,WX4880,WX4542);
  nand NAND2_2485(II14283,WX4880,II14282);
  nand NAND2_2486(II14284,WX4542,II14282);
  nand NAND2_2487(II14281,II14283,II14284);
  nand NAND2_2488(II14289,WX4606,II14281);
  nand NAND2_2489(II14290,WX4606,II14289);
  nand NAND2_2490(II14291,II14281,II14289);
  nand NAND2_2491(II14280,II14290,II14291);
  nand NAND2_2492(II14297,WX4670,WX4734);
  nand NAND2_2493(II14298,WX4670,II14297);
  nand NAND2_2494(II14299,WX4734,II14297);
  nand NAND2_2495(II14296,II14298,II14299);
  nand NAND2_2496(II14304,II14280,II14296);
  nand NAND2_2497(II14305,II14280,II14304);
  nand NAND2_2498(II14306,II14296,II14304);
  nand NAND2_2499(WX4788,II14305,II14306);
  nand NAND2_2500(II14313,WX4880,WX4544);
  nand NAND2_2501(II14314,WX4880,II14313);
  nand NAND2_2502(II14315,WX4544,II14313);
  nand NAND2_2503(II14312,II14314,II14315);
  nand NAND2_2504(II14320,WX4608,II14312);
  nand NAND2_2505(II14321,WX4608,II14320);
  nand NAND2_2506(II14322,II14312,II14320);
  nand NAND2_2507(II14311,II14321,II14322);
  nand NAND2_2508(II14328,WX4672,WX4736);
  nand NAND2_2509(II14329,WX4672,II14328);
  nand NAND2_2510(II14330,WX4736,II14328);
  nand NAND2_2511(II14327,II14329,II14330);
  nand NAND2_2512(II14335,II14311,II14327);
  nand NAND2_2513(II14336,II14311,II14335);
  nand NAND2_2514(II14337,II14327,II14335);
  nand NAND2_2515(WX4789,II14336,II14337);
  nand NAND2_2516(II14344,WX4880,WX4546);
  nand NAND2_2517(II14345,WX4880,II14344);
  nand NAND2_2518(II14346,WX4546,II14344);
  nand NAND2_2519(II14343,II14345,II14346);
  nand NAND2_2520(II14351,WX4610,II14343);
  nand NAND2_2521(II14352,WX4610,II14351);
  nand NAND2_2522(II14353,II14343,II14351);
  nand NAND2_2523(II14342,II14352,II14353);
  nand NAND2_2524(II14359,WX4674,WX4738);
  nand NAND2_2525(II14360,WX4674,II14359);
  nand NAND2_2526(II14361,WX4738,II14359);
  nand NAND2_2527(II14358,II14360,II14361);
  nand NAND2_2528(II14366,II14342,II14358);
  nand NAND2_2529(II14367,II14342,II14366);
  nand NAND2_2530(II14368,II14358,II14366);
  nand NAND2_2531(WX4790,II14367,II14368);
  nand NAND2_2532(II14375,WX4880,WX4548);
  nand NAND2_2533(II14376,WX4880,II14375);
  nand NAND2_2534(II14377,WX4548,II14375);
  nand NAND2_2535(II14374,II14376,II14377);
  nand NAND2_2536(II14382,WX4612,II14374);
  nand NAND2_2537(II14383,WX4612,II14382);
  nand NAND2_2538(II14384,II14374,II14382);
  nand NAND2_2539(II14373,II14383,II14384);
  nand NAND2_2540(II14390,WX4676,WX4740);
  nand NAND2_2541(II14391,WX4676,II14390);
  nand NAND2_2542(II14392,WX4740,II14390);
  nand NAND2_2543(II14389,II14391,II14392);
  nand NAND2_2544(II14397,II14373,II14389);
  nand NAND2_2545(II14398,II14373,II14397);
  nand NAND2_2546(II14399,II14389,II14397);
  nand NAND2_2547(WX4791,II14398,II14399);
  nand NAND2_2548(II14406,WX4880,WX4550);
  nand NAND2_2549(II14407,WX4880,II14406);
  nand NAND2_2550(II14408,WX4550,II14406);
  nand NAND2_2551(II14405,II14407,II14408);
  nand NAND2_2552(II14413,WX4614,II14405);
  nand NAND2_2553(II14414,WX4614,II14413);
  nand NAND2_2554(II14415,II14405,II14413);
  nand NAND2_2555(II14404,II14414,II14415);
  nand NAND2_2556(II14421,WX4678,WX4742);
  nand NAND2_2557(II14422,WX4678,II14421);
  nand NAND2_2558(II14423,WX4742,II14421);
  nand NAND2_2559(II14420,II14422,II14423);
  nand NAND2_2560(II14428,II14404,II14420);
  nand NAND2_2561(II14429,II14404,II14428);
  nand NAND2_2562(II14430,II14420,II14428);
  nand NAND2_2563(WX4792,II14429,II14430);
  nand NAND2_2564(II14437,WX4880,WX4552);
  nand NAND2_2565(II14438,WX4880,II14437);
  nand NAND2_2566(II14439,WX4552,II14437);
  nand NAND2_2567(II14436,II14438,II14439);
  nand NAND2_2568(II14444,WX4616,II14436);
  nand NAND2_2569(II14445,WX4616,II14444);
  nand NAND2_2570(II14446,II14436,II14444);
  nand NAND2_2571(II14435,II14445,II14446);
  nand NAND2_2572(II14452,WX4680,WX4744);
  nand NAND2_2573(II14453,WX4680,II14452);
  nand NAND2_2574(II14454,WX4744,II14452);
  nand NAND2_2575(II14451,II14453,II14454);
  nand NAND2_2576(II14459,II14435,II14451);
  nand NAND2_2577(II14460,II14435,II14459);
  nand NAND2_2578(II14461,II14451,II14459);
  nand NAND2_2579(WX4793,II14460,II14461);
  nand NAND2_2580(II14468,WX4880,WX4554);
  nand NAND2_2581(II14469,WX4880,II14468);
  nand NAND2_2582(II14470,WX4554,II14468);
  nand NAND2_2583(II14467,II14469,II14470);
  nand NAND2_2584(II14475,WX4618,II14467);
  nand NAND2_2585(II14476,WX4618,II14475);
  nand NAND2_2586(II14477,II14467,II14475);
  nand NAND2_2587(II14466,II14476,II14477);
  nand NAND2_2588(II14483,WX4682,WX4746);
  nand NAND2_2589(II14484,WX4682,II14483);
  nand NAND2_2590(II14485,WX4746,II14483);
  nand NAND2_2591(II14482,II14484,II14485);
  nand NAND2_2592(II14490,II14466,II14482);
  nand NAND2_2593(II14491,II14466,II14490);
  nand NAND2_2594(II14492,II14482,II14490);
  nand NAND2_2595(WX4794,II14491,II14492);
  nand NAND2_2596(II14499,WX4881,WX4556);
  nand NAND2_2597(II14500,WX4881,II14499);
  nand NAND2_2598(II14501,WX4556,II14499);
  nand NAND2_2599(II14498,II14500,II14501);
  nand NAND2_2600(II14506,WX4620,II14498);
  nand NAND2_2601(II14507,WX4620,II14506);
  nand NAND2_2602(II14508,II14498,II14506);
  nand NAND2_2603(II14497,II14507,II14508);
  nand NAND2_2604(II14514,WX4684,WX4748);
  nand NAND2_2605(II14515,WX4684,II14514);
  nand NAND2_2606(II14516,WX4748,II14514);
  nand NAND2_2607(II14513,II14515,II14516);
  nand NAND2_2608(II14521,II14497,II14513);
  nand NAND2_2609(II14522,II14497,II14521);
  nand NAND2_2610(II14523,II14513,II14521);
  nand NAND2_2611(WX4795,II14522,II14523);
  nand NAND2_2612(II14530,WX4881,WX4558);
  nand NAND2_2613(II14531,WX4881,II14530);
  nand NAND2_2614(II14532,WX4558,II14530);
  nand NAND2_2615(II14529,II14531,II14532);
  nand NAND2_2616(II14537,WX4622,II14529);
  nand NAND2_2617(II14538,WX4622,II14537);
  nand NAND2_2618(II14539,II14529,II14537);
  nand NAND2_2619(II14528,II14538,II14539);
  nand NAND2_2620(II14545,WX4686,WX4750);
  nand NAND2_2621(II14546,WX4686,II14545);
  nand NAND2_2622(II14547,WX4750,II14545);
  nand NAND2_2623(II14544,II14546,II14547);
  nand NAND2_2624(II14552,II14528,II14544);
  nand NAND2_2625(II14553,II14528,II14552);
  nand NAND2_2626(II14554,II14544,II14552);
  nand NAND2_2627(WX4796,II14553,II14554);
  nand NAND2_2628(II14561,WX4881,WX4560);
  nand NAND2_2629(II14562,WX4881,II14561);
  nand NAND2_2630(II14563,WX4560,II14561);
  nand NAND2_2631(II14560,II14562,II14563);
  nand NAND2_2632(II14568,WX4624,II14560);
  nand NAND2_2633(II14569,WX4624,II14568);
  nand NAND2_2634(II14570,II14560,II14568);
  nand NAND2_2635(II14559,II14569,II14570);
  nand NAND2_2636(II14576,WX4688,WX4752);
  nand NAND2_2637(II14577,WX4688,II14576);
  nand NAND2_2638(II14578,WX4752,II14576);
  nand NAND2_2639(II14575,II14577,II14578);
  nand NAND2_2640(II14583,II14559,II14575);
  nand NAND2_2641(II14584,II14559,II14583);
  nand NAND2_2642(II14585,II14575,II14583);
  nand NAND2_2643(WX4797,II14584,II14585);
  nand NAND2_2644(II14592,WX4881,WX4562);
  nand NAND2_2645(II14593,WX4881,II14592);
  nand NAND2_2646(II14594,WX4562,II14592);
  nand NAND2_2647(II14591,II14593,II14594);
  nand NAND2_2648(II14599,WX4626,II14591);
  nand NAND2_2649(II14600,WX4626,II14599);
  nand NAND2_2650(II14601,II14591,II14599);
  nand NAND2_2651(II14590,II14600,II14601);
  nand NAND2_2652(II14607,WX4690,WX4754);
  nand NAND2_2653(II14608,WX4690,II14607);
  nand NAND2_2654(II14609,WX4754,II14607);
  nand NAND2_2655(II14606,II14608,II14609);
  nand NAND2_2656(II14614,II14590,II14606);
  nand NAND2_2657(II14615,II14590,II14614);
  nand NAND2_2658(II14616,II14606,II14614);
  nand NAND2_2659(WX4798,II14615,II14616);
  nand NAND2_2660(II14623,WX4881,WX4564);
  nand NAND2_2661(II14624,WX4881,II14623);
  nand NAND2_2662(II14625,WX4564,II14623);
  nand NAND2_2663(II14622,II14624,II14625);
  nand NAND2_2664(II14630,WX4628,II14622);
  nand NAND2_2665(II14631,WX4628,II14630);
  nand NAND2_2666(II14632,II14622,II14630);
  nand NAND2_2667(II14621,II14631,II14632);
  nand NAND2_2668(II14638,WX4692,WX4756);
  nand NAND2_2669(II14639,WX4692,II14638);
  nand NAND2_2670(II14640,WX4756,II14638);
  nand NAND2_2671(II14637,II14639,II14640);
  nand NAND2_2672(II14645,II14621,II14637);
  nand NAND2_2673(II14646,II14621,II14645);
  nand NAND2_2674(II14647,II14637,II14645);
  nand NAND2_2675(WX4799,II14646,II14647);
  nand NAND2_2676(II14654,WX4881,WX4566);
  nand NAND2_2677(II14655,WX4881,II14654);
  nand NAND2_2678(II14656,WX4566,II14654);
  nand NAND2_2679(II14653,II14655,II14656);
  nand NAND2_2680(II14661,WX4630,II14653);
  nand NAND2_2681(II14662,WX4630,II14661);
  nand NAND2_2682(II14663,II14653,II14661);
  nand NAND2_2683(II14652,II14662,II14663);
  nand NAND2_2684(II14669,WX4694,WX4758);
  nand NAND2_2685(II14670,WX4694,II14669);
  nand NAND2_2686(II14671,WX4758,II14669);
  nand NAND2_2687(II14668,II14670,II14671);
  nand NAND2_2688(II14676,II14652,II14668);
  nand NAND2_2689(II14677,II14652,II14676);
  nand NAND2_2690(II14678,II14668,II14676);
  nand NAND2_2691(WX4800,II14677,II14678);
  nand NAND2_2692(II14685,WX4881,WX4568);
  nand NAND2_2693(II14686,WX4881,II14685);
  nand NAND2_2694(II14687,WX4568,II14685);
  nand NAND2_2695(II14684,II14686,II14687);
  nand NAND2_2696(II14692,WX4632,II14684);
  nand NAND2_2697(II14693,WX4632,II14692);
  nand NAND2_2698(II14694,II14684,II14692);
  nand NAND2_2699(II14683,II14693,II14694);
  nand NAND2_2700(II14700,WX4696,WX4760);
  nand NAND2_2701(II14701,WX4696,II14700);
  nand NAND2_2702(II14702,WX4760,II14700);
  nand NAND2_2703(II14699,II14701,II14702);
  nand NAND2_2704(II14707,II14683,II14699);
  nand NAND2_2705(II14708,II14683,II14707);
  nand NAND2_2706(II14709,II14699,II14707);
  nand NAND2_2707(WX4801,II14708,II14709);
  nand NAND2_2708(II14716,WX4881,WX4570);
  nand NAND2_2709(II14717,WX4881,II14716);
  nand NAND2_2710(II14718,WX4570,II14716);
  nand NAND2_2711(II14715,II14717,II14718);
  nand NAND2_2712(II14723,WX4634,II14715);
  nand NAND2_2713(II14724,WX4634,II14723);
  nand NAND2_2714(II14725,II14715,II14723);
  nand NAND2_2715(II14714,II14724,II14725);
  nand NAND2_2716(II14731,WX4698,WX4762);
  nand NAND2_2717(II14732,WX4698,II14731);
  nand NAND2_2718(II14733,WX4762,II14731);
  nand NAND2_2719(II14730,II14732,II14733);
  nand NAND2_2720(II14738,II14714,II14730);
  nand NAND2_2721(II14739,II14714,II14738);
  nand NAND2_2722(II14740,II14730,II14738);
  nand NAND2_2723(WX4802,II14739,II14740);
  nand NAND2_2724(II14747,WX4881,WX4572);
  nand NAND2_2725(II14748,WX4881,II14747);
  nand NAND2_2726(II14749,WX4572,II14747);
  nand NAND2_2727(II14746,II14748,II14749);
  nand NAND2_2728(II14754,WX4636,II14746);
  nand NAND2_2729(II14755,WX4636,II14754);
  nand NAND2_2730(II14756,II14746,II14754);
  nand NAND2_2731(II14745,II14755,II14756);
  nand NAND2_2732(II14762,WX4700,WX4764);
  nand NAND2_2733(II14763,WX4700,II14762);
  nand NAND2_2734(II14764,WX4764,II14762);
  nand NAND2_2735(II14761,II14763,II14764);
  nand NAND2_2736(II14769,II14745,II14761);
  nand NAND2_2737(II14770,II14745,II14769);
  nand NAND2_2738(II14771,II14761,II14769);
  nand NAND2_2739(WX4803,II14770,II14771);
  nand NAND2_2740(II14778,WX4881,WX4574);
  nand NAND2_2741(II14779,WX4881,II14778);
  nand NAND2_2742(II14780,WX4574,II14778);
  nand NAND2_2743(II14777,II14779,II14780);
  nand NAND2_2744(II14785,WX4638,II14777);
  nand NAND2_2745(II14786,WX4638,II14785);
  nand NAND2_2746(II14787,II14777,II14785);
  nand NAND2_2747(II14776,II14786,II14787);
  nand NAND2_2748(II14793,WX4702,WX4766);
  nand NAND2_2749(II14794,WX4702,II14793);
  nand NAND2_2750(II14795,WX4766,II14793);
  nand NAND2_2751(II14792,II14794,II14795);
  nand NAND2_2752(II14800,II14776,II14792);
  nand NAND2_2753(II14801,II14776,II14800);
  nand NAND2_2754(II14802,II14792,II14800);
  nand NAND2_2755(WX4804,II14801,II14802);
  nand NAND2_2756(II14809,WX4881,WX4576);
  nand NAND2_2757(II14810,WX4881,II14809);
  nand NAND2_2758(II14811,WX4576,II14809);
  nand NAND2_2759(II14808,II14810,II14811);
  nand NAND2_2760(II14816,WX4640,II14808);
  nand NAND2_2761(II14817,WX4640,II14816);
  nand NAND2_2762(II14818,II14808,II14816);
  nand NAND2_2763(II14807,II14817,II14818);
  nand NAND2_2764(II14824,WX4704,WX4768);
  nand NAND2_2765(II14825,WX4704,II14824);
  nand NAND2_2766(II14826,WX4768,II14824);
  nand NAND2_2767(II14823,II14825,II14826);
  nand NAND2_2768(II14831,II14807,II14823);
  nand NAND2_2769(II14832,II14807,II14831);
  nand NAND2_2770(II14833,II14823,II14831);
  nand NAND2_2771(WX4805,II14832,II14833);
  nand NAND2_2772(II14840,WX4881,WX4578);
  nand NAND2_2773(II14841,WX4881,II14840);
  nand NAND2_2774(II14842,WX4578,II14840);
  nand NAND2_2775(II14839,II14841,II14842);
  nand NAND2_2776(II14847,WX4642,II14839);
  nand NAND2_2777(II14848,WX4642,II14847);
  nand NAND2_2778(II14849,II14839,II14847);
  nand NAND2_2779(II14838,II14848,II14849);
  nand NAND2_2780(II14855,WX4706,WX4770);
  nand NAND2_2781(II14856,WX4706,II14855);
  nand NAND2_2782(II14857,WX4770,II14855);
  nand NAND2_2783(II14854,II14856,II14857);
  nand NAND2_2784(II14862,II14838,II14854);
  nand NAND2_2785(II14863,II14838,II14862);
  nand NAND2_2786(II14864,II14854,II14862);
  nand NAND2_2787(WX4806,II14863,II14864);
  nand NAND2_2788(II14871,WX4881,WX4580);
  nand NAND2_2789(II14872,WX4881,II14871);
  nand NAND2_2790(II14873,WX4580,II14871);
  nand NAND2_2791(II14870,II14872,II14873);
  nand NAND2_2792(II14878,WX4644,II14870);
  nand NAND2_2793(II14879,WX4644,II14878);
  nand NAND2_2794(II14880,II14870,II14878);
  nand NAND2_2795(II14869,II14879,II14880);
  nand NAND2_2796(II14886,WX4708,WX4772);
  nand NAND2_2797(II14887,WX4708,II14886);
  nand NAND2_2798(II14888,WX4772,II14886);
  nand NAND2_2799(II14885,II14887,II14888);
  nand NAND2_2800(II14893,II14869,II14885);
  nand NAND2_2801(II14894,II14869,II14893);
  nand NAND2_2802(II14895,II14885,II14893);
  nand NAND2_2803(WX4807,II14894,II14895);
  nand NAND2_2804(II14902,WX4881,WX4582);
  nand NAND2_2805(II14903,WX4881,II14902);
  nand NAND2_2806(II14904,WX4582,II14902);
  nand NAND2_2807(II14901,II14903,II14904);
  nand NAND2_2808(II14909,WX4646,II14901);
  nand NAND2_2809(II14910,WX4646,II14909);
  nand NAND2_2810(II14911,II14901,II14909);
  nand NAND2_2811(II14900,II14910,II14911);
  nand NAND2_2812(II14917,WX4710,WX4774);
  nand NAND2_2813(II14918,WX4710,II14917);
  nand NAND2_2814(II14919,WX4774,II14917);
  nand NAND2_2815(II14916,II14918,II14919);
  nand NAND2_2816(II14924,II14900,II14916);
  nand NAND2_2817(II14925,II14900,II14924);
  nand NAND2_2818(II14926,II14916,II14924);
  nand NAND2_2819(WX4808,II14925,II14926);
  nand NAND2_2820(II14933,WX4881,WX4584);
  nand NAND2_2821(II14934,WX4881,II14933);
  nand NAND2_2822(II14935,WX4584,II14933);
  nand NAND2_2823(II14932,II14934,II14935);
  nand NAND2_2824(II14940,WX4648,II14932);
  nand NAND2_2825(II14941,WX4648,II14940);
  nand NAND2_2826(II14942,II14932,II14940);
  nand NAND2_2827(II14931,II14941,II14942);
  nand NAND2_2828(II14948,WX4712,WX4776);
  nand NAND2_2829(II14949,WX4712,II14948);
  nand NAND2_2830(II14950,WX4776,II14948);
  nand NAND2_2831(II14947,II14949,II14950);
  nand NAND2_2832(II14955,II14931,II14947);
  nand NAND2_2833(II14956,II14931,II14955);
  nand NAND2_2834(II14957,II14947,II14955);
  nand NAND2_2835(WX4809,II14956,II14957);
  nand NAND2_2836(II14964,WX4881,WX4586);
  nand NAND2_2837(II14965,WX4881,II14964);
  nand NAND2_2838(II14966,WX4586,II14964);
  nand NAND2_2839(II14963,II14965,II14966);
  nand NAND2_2840(II14971,WX4650,II14963);
  nand NAND2_2841(II14972,WX4650,II14971);
  nand NAND2_2842(II14973,II14963,II14971);
  nand NAND2_2843(II14962,II14972,II14973);
  nand NAND2_2844(II14979,WX4714,WX4778);
  nand NAND2_2845(II14980,WX4714,II14979);
  nand NAND2_2846(II14981,WX4778,II14979);
  nand NAND2_2847(II14978,II14980,II14981);
  nand NAND2_2848(II14986,II14962,II14978);
  nand NAND2_2849(II14987,II14962,II14986);
  nand NAND2_2850(II14988,II14978,II14986);
  nand NAND2_2851(WX4810,II14987,II14988);
  nand NAND2_2852(II15067,WX4459,WX4364);
  nand NAND2_2853(II15068,WX4459,II15067);
  nand NAND2_2854(II15069,WX4364,II15067);
  nand NAND2_2855(WX4885,II15068,II15069);
  nand NAND2_2856(II15080,WX4460,WX4366);
  nand NAND2_2857(II15081,WX4460,II15080);
  nand NAND2_2858(II15082,WX4366,II15080);
  nand NAND2_2859(WX4892,II15081,II15082);
  nand NAND2_2860(II15093,WX4461,WX4368);
  nand NAND2_2861(II15094,WX4461,II15093);
  nand NAND2_2862(II15095,WX4368,II15093);
  nand NAND2_2863(WX4899,II15094,II15095);
  nand NAND2_2864(II15106,WX4462,WX4370);
  nand NAND2_2865(II15107,WX4462,II15106);
  nand NAND2_2866(II15108,WX4370,II15106);
  nand NAND2_2867(WX4906,II15107,II15108);
  nand NAND2_2868(II15119,WX4463,WX4372);
  nand NAND2_2869(II15120,WX4463,II15119);
  nand NAND2_2870(II15121,WX4372,II15119);
  nand NAND2_2871(WX4913,II15120,II15121);
  nand NAND2_2872(II15132,WX4464,WX4374);
  nand NAND2_2873(II15133,WX4464,II15132);
  nand NAND2_2874(II15134,WX4374,II15132);
  nand NAND2_2875(WX4920,II15133,II15134);
  nand NAND2_2876(II15145,WX4465,WX4376);
  nand NAND2_2877(II15146,WX4465,II15145);
  nand NAND2_2878(II15147,WX4376,II15145);
  nand NAND2_2879(WX4927,II15146,II15147);
  nand NAND2_2880(II15158,WX4466,WX4378);
  nand NAND2_2881(II15159,WX4466,II15158);
  nand NAND2_2882(II15160,WX4378,II15158);
  nand NAND2_2883(WX4934,II15159,II15160);
  nand NAND2_2884(II15171,WX4467,WX4380);
  nand NAND2_2885(II15172,WX4467,II15171);
  nand NAND2_2886(II15173,WX4380,II15171);
  nand NAND2_2887(WX4941,II15172,II15173);
  nand NAND2_2888(II15184,WX4468,WX4382);
  nand NAND2_2889(II15185,WX4468,II15184);
  nand NAND2_2890(II15186,WX4382,II15184);
  nand NAND2_2891(WX4948,II15185,II15186);
  nand NAND2_2892(II15197,WX4469,WX4384);
  nand NAND2_2893(II15198,WX4469,II15197);
  nand NAND2_2894(II15199,WX4384,II15197);
  nand NAND2_2895(WX4955,II15198,II15199);
  nand NAND2_2896(II15210,WX4470,WX4386);
  nand NAND2_2897(II15211,WX4470,II15210);
  nand NAND2_2898(II15212,WX4386,II15210);
  nand NAND2_2899(WX4962,II15211,II15212);
  nand NAND2_2900(II15223,WX4471,WX4388);
  nand NAND2_2901(II15224,WX4471,II15223);
  nand NAND2_2902(II15225,WX4388,II15223);
  nand NAND2_2903(WX4969,II15224,II15225);
  nand NAND2_2904(II15236,WX4472,WX4390);
  nand NAND2_2905(II15237,WX4472,II15236);
  nand NAND2_2906(II15238,WX4390,II15236);
  nand NAND2_2907(WX4976,II15237,II15238);
  nand NAND2_2908(II15249,WX4473,WX4392);
  nand NAND2_2909(II15250,WX4473,II15249);
  nand NAND2_2910(II15251,WX4392,II15249);
  nand NAND2_2911(WX4983,II15250,II15251);
  nand NAND2_2912(II15262,WX4474,WX4394);
  nand NAND2_2913(II15263,WX4474,II15262);
  nand NAND2_2914(II15264,WX4394,II15262);
  nand NAND2_2915(WX4990,II15263,II15264);
  nand NAND2_2916(II15275,WX4475,WX4396);
  nand NAND2_2917(II15276,WX4475,II15275);
  nand NAND2_2918(II15277,WX4396,II15275);
  nand NAND2_2919(WX4997,II15276,II15277);
  nand NAND2_2920(II15288,WX4476,WX4398);
  nand NAND2_2921(II15289,WX4476,II15288);
  nand NAND2_2922(II15290,WX4398,II15288);
  nand NAND2_2923(WX5004,II15289,II15290);
  nand NAND2_2924(II15301,WX4477,WX4400);
  nand NAND2_2925(II15302,WX4477,II15301);
  nand NAND2_2926(II15303,WX4400,II15301);
  nand NAND2_2927(WX5011,II15302,II15303);
  nand NAND2_2928(II15314,WX4478,WX4402);
  nand NAND2_2929(II15315,WX4478,II15314);
  nand NAND2_2930(II15316,WX4402,II15314);
  nand NAND2_2931(WX5018,II15315,II15316);
  nand NAND2_2932(II15327,WX4479,WX4404);
  nand NAND2_2933(II15328,WX4479,II15327);
  nand NAND2_2934(II15329,WX4404,II15327);
  nand NAND2_2935(WX5025,II15328,II15329);
  nand NAND2_2936(II15340,WX4480,WX4406);
  nand NAND2_2937(II15341,WX4480,II15340);
  nand NAND2_2938(II15342,WX4406,II15340);
  nand NAND2_2939(WX5032,II15341,II15342);
  nand NAND2_2940(II15353,WX4481,WX4408);
  nand NAND2_2941(II15354,WX4481,II15353);
  nand NAND2_2942(II15355,WX4408,II15353);
  nand NAND2_2943(WX5039,II15354,II15355);
  nand NAND2_2944(II15366,WX4482,WX4410);
  nand NAND2_2945(II15367,WX4482,II15366);
  nand NAND2_2946(II15368,WX4410,II15366);
  nand NAND2_2947(WX5046,II15367,II15368);
  nand NAND2_2948(II15379,WX4483,WX4412);
  nand NAND2_2949(II15380,WX4483,II15379);
  nand NAND2_2950(II15381,WX4412,II15379);
  nand NAND2_2951(WX5053,II15380,II15381);
  nand NAND2_2952(II15392,WX4484,WX4414);
  nand NAND2_2953(II15393,WX4484,II15392);
  nand NAND2_2954(II15394,WX4414,II15392);
  nand NAND2_2955(WX5060,II15393,II15394);
  nand NAND2_2956(II15405,WX4485,WX4416);
  nand NAND2_2957(II15406,WX4485,II15405);
  nand NAND2_2958(II15407,WX4416,II15405);
  nand NAND2_2959(WX5067,II15406,II15407);
  nand NAND2_2960(II15418,WX4486,WX4418);
  nand NAND2_2961(II15419,WX4486,II15418);
  nand NAND2_2962(II15420,WX4418,II15418);
  nand NAND2_2963(WX5074,II15419,II15420);
  nand NAND2_2964(II15431,WX4487,WX4420);
  nand NAND2_2965(II15432,WX4487,II15431);
  nand NAND2_2966(II15433,WX4420,II15431);
  nand NAND2_2967(WX5081,II15432,II15433);
  nand NAND2_2968(II15444,WX4488,WX4422);
  nand NAND2_2969(II15445,WX4488,II15444);
  nand NAND2_2970(II15446,WX4422,II15444);
  nand NAND2_2971(WX5088,II15445,II15446);
  nand NAND2_2972(II15457,WX4489,WX4424);
  nand NAND2_2973(II15458,WX4489,II15457);
  nand NAND2_2974(II15459,WX4424,II15457);
  nand NAND2_2975(WX5095,II15458,II15459);
  nand NAND2_2976(II15470,WX4490,WX4426);
  nand NAND2_2977(II15471,WX4490,II15470);
  nand NAND2_2978(II15472,WX4426,II15470);
  nand NAND2_2979(WX5102,II15471,II15472);
  nand NAND2_2980(II15485,WX4506,CRC_OUT_6_31);
  nand NAND2_2981(II15486,WX4506,II15485);
  nand NAND2_2982(II15487,CRC_OUT_6_31,II15485);
  nand NAND2_2983(II15484,II15486,II15487);
  nand NAND2_2984(II15492,CRC_OUT_6_15,II15484);
  nand NAND2_2985(II15493,CRC_OUT_6_15,II15492);
  nand NAND2_2986(II15494,II15484,II15492);
  nand NAND2_2987(WX5110,II15493,II15494);
  nand NAND2_2988(II15500,WX4511,CRC_OUT_6_31);
  nand NAND2_2989(II15501,WX4511,II15500);
  nand NAND2_2990(II15502,CRC_OUT_6_31,II15500);
  nand NAND2_2991(II15499,II15501,II15502);
  nand NAND2_2992(II15507,CRC_OUT_6_10,II15499);
  nand NAND2_2993(II15508,CRC_OUT_6_10,II15507);
  nand NAND2_2994(II15509,II15499,II15507);
  nand NAND2_2995(WX5111,II15508,II15509);
  nand NAND2_2996(II15515,WX4518,CRC_OUT_6_31);
  nand NAND2_2997(II15516,WX4518,II15515);
  nand NAND2_2998(II15517,CRC_OUT_6_31,II15515);
  nand NAND2_2999(II15514,II15516,II15517);
  nand NAND2_3000(II15522,CRC_OUT_6_3,II15514);
  nand NAND2_3001(II15523,CRC_OUT_6_3,II15522);
  nand NAND2_3002(II15524,II15514,II15522);
  nand NAND2_3003(WX5112,II15523,II15524);
  nand NAND2_3004(II15529,WX4522,CRC_OUT_6_31);
  nand NAND2_3005(II15530,WX4522,II15529);
  nand NAND2_3006(II15531,CRC_OUT_6_31,II15529);
  nand NAND2_3007(WX5113,II15530,II15531);
  nand NAND2_3008(II15536,WX4491,CRC_OUT_6_30);
  nand NAND2_3009(II15537,WX4491,II15536);
  nand NAND2_3010(II15538,CRC_OUT_6_30,II15536);
  nand NAND2_3011(WX5114,II15537,II15538);
  nand NAND2_3012(II15543,WX4492,CRC_OUT_6_29);
  nand NAND2_3013(II15544,WX4492,II15543);
  nand NAND2_3014(II15545,CRC_OUT_6_29,II15543);
  nand NAND2_3015(WX5115,II15544,II15545);
  nand NAND2_3016(II15550,WX4493,CRC_OUT_6_28);
  nand NAND2_3017(II15551,WX4493,II15550);
  nand NAND2_3018(II15552,CRC_OUT_6_28,II15550);
  nand NAND2_3019(WX5116,II15551,II15552);
  nand NAND2_3020(II15557,WX4494,CRC_OUT_6_27);
  nand NAND2_3021(II15558,WX4494,II15557);
  nand NAND2_3022(II15559,CRC_OUT_6_27,II15557);
  nand NAND2_3023(WX5117,II15558,II15559);
  nand NAND2_3024(II15564,WX4495,CRC_OUT_6_26);
  nand NAND2_3025(II15565,WX4495,II15564);
  nand NAND2_3026(II15566,CRC_OUT_6_26,II15564);
  nand NAND2_3027(WX5118,II15565,II15566);
  nand NAND2_3028(II15571,WX4496,CRC_OUT_6_25);
  nand NAND2_3029(II15572,WX4496,II15571);
  nand NAND2_3030(II15573,CRC_OUT_6_25,II15571);
  nand NAND2_3031(WX5119,II15572,II15573);
  nand NAND2_3032(II15578,WX4497,CRC_OUT_6_24);
  nand NAND2_3033(II15579,WX4497,II15578);
  nand NAND2_3034(II15580,CRC_OUT_6_24,II15578);
  nand NAND2_3035(WX5120,II15579,II15580);
  nand NAND2_3036(II15585,WX4498,CRC_OUT_6_23);
  nand NAND2_3037(II15586,WX4498,II15585);
  nand NAND2_3038(II15587,CRC_OUT_6_23,II15585);
  nand NAND2_3039(WX5121,II15586,II15587);
  nand NAND2_3040(II15592,WX4499,CRC_OUT_6_22);
  nand NAND2_3041(II15593,WX4499,II15592);
  nand NAND2_3042(II15594,CRC_OUT_6_22,II15592);
  nand NAND2_3043(WX5122,II15593,II15594);
  nand NAND2_3044(II15599,WX4500,CRC_OUT_6_21);
  nand NAND2_3045(II15600,WX4500,II15599);
  nand NAND2_3046(II15601,CRC_OUT_6_21,II15599);
  nand NAND2_3047(WX5123,II15600,II15601);
  nand NAND2_3048(II15606,WX4501,CRC_OUT_6_20);
  nand NAND2_3049(II15607,WX4501,II15606);
  nand NAND2_3050(II15608,CRC_OUT_6_20,II15606);
  nand NAND2_3051(WX5124,II15607,II15608);
  nand NAND2_3052(II15613,WX4502,CRC_OUT_6_19);
  nand NAND2_3053(II15614,WX4502,II15613);
  nand NAND2_3054(II15615,CRC_OUT_6_19,II15613);
  nand NAND2_3055(WX5125,II15614,II15615);
  nand NAND2_3056(II15620,WX4503,CRC_OUT_6_18);
  nand NAND2_3057(II15621,WX4503,II15620);
  nand NAND2_3058(II15622,CRC_OUT_6_18,II15620);
  nand NAND2_3059(WX5126,II15621,II15622);
  nand NAND2_3060(II15627,WX4504,CRC_OUT_6_17);
  nand NAND2_3061(II15628,WX4504,II15627);
  nand NAND2_3062(II15629,CRC_OUT_6_17,II15627);
  nand NAND2_3063(WX5127,II15628,II15629);
  nand NAND2_3064(II15634,WX4505,CRC_OUT_6_16);
  nand NAND2_3065(II15635,WX4505,II15634);
  nand NAND2_3066(II15636,CRC_OUT_6_16,II15634);
  nand NAND2_3067(WX5128,II15635,II15636);
  nand NAND2_3068(II15641,WX4507,CRC_OUT_6_14);
  nand NAND2_3069(II15642,WX4507,II15641);
  nand NAND2_3070(II15643,CRC_OUT_6_14,II15641);
  nand NAND2_3071(WX5129,II15642,II15643);
  nand NAND2_3072(II15648,WX4508,CRC_OUT_6_13);
  nand NAND2_3073(II15649,WX4508,II15648);
  nand NAND2_3074(II15650,CRC_OUT_6_13,II15648);
  nand NAND2_3075(WX5130,II15649,II15650);
  nand NAND2_3076(II15655,WX4509,CRC_OUT_6_12);
  nand NAND2_3077(II15656,WX4509,II15655);
  nand NAND2_3078(II15657,CRC_OUT_6_12,II15655);
  nand NAND2_3079(WX5131,II15656,II15657);
  nand NAND2_3080(II15662,WX4510,CRC_OUT_6_11);
  nand NAND2_3081(II15663,WX4510,II15662);
  nand NAND2_3082(II15664,CRC_OUT_6_11,II15662);
  nand NAND2_3083(WX5132,II15663,II15664);
  nand NAND2_3084(II15669,WX4512,CRC_OUT_6_9);
  nand NAND2_3085(II15670,WX4512,II15669);
  nand NAND2_3086(II15671,CRC_OUT_6_9,II15669);
  nand NAND2_3087(WX5133,II15670,II15671);
  nand NAND2_3088(II15676,WX4513,CRC_OUT_6_8);
  nand NAND2_3089(II15677,WX4513,II15676);
  nand NAND2_3090(II15678,CRC_OUT_6_8,II15676);
  nand NAND2_3091(WX5134,II15677,II15678);
  nand NAND2_3092(II15683,WX4514,CRC_OUT_6_7);
  nand NAND2_3093(II15684,WX4514,II15683);
  nand NAND2_3094(II15685,CRC_OUT_6_7,II15683);
  nand NAND2_3095(WX5135,II15684,II15685);
  nand NAND2_3096(II15690,WX4515,CRC_OUT_6_6);
  nand NAND2_3097(II15691,WX4515,II15690);
  nand NAND2_3098(II15692,CRC_OUT_6_6,II15690);
  nand NAND2_3099(WX5136,II15691,II15692);
  nand NAND2_3100(II15697,WX4516,CRC_OUT_6_5);
  nand NAND2_3101(II15698,WX4516,II15697);
  nand NAND2_3102(II15699,CRC_OUT_6_5,II15697);
  nand NAND2_3103(WX5137,II15698,II15699);
  nand NAND2_3104(II15704,WX4517,CRC_OUT_6_4);
  nand NAND2_3105(II15705,WX4517,II15704);
  nand NAND2_3106(II15706,CRC_OUT_6_4,II15704);
  nand NAND2_3107(WX5138,II15705,II15706);
  nand NAND2_3108(II15711,WX4519,CRC_OUT_6_2);
  nand NAND2_3109(II15712,WX4519,II15711);
  nand NAND2_3110(II15713,CRC_OUT_6_2,II15711);
  nand NAND2_3111(WX5139,II15712,II15713);
  nand NAND2_3112(II15718,WX4520,CRC_OUT_6_1);
  nand NAND2_3113(II15719,WX4520,II15718);
  nand NAND2_3114(II15720,CRC_OUT_6_1,II15718);
  nand NAND2_3115(WX5140,II15719,II15720);
  nand NAND2_3116(II15725,WX4521,CRC_OUT_6_0);
  nand NAND2_3117(II15726,WX4521,II15725);
  nand NAND2_3118(II15727,CRC_OUT_6_0,II15725);
  nand NAND2_3119(WX5141,II15726,II15727);
  nand NAND2_3120(II18008,WX6173,WX5817);
  nand NAND2_3121(II18009,WX6173,II18008);
  nand NAND2_3122(II18010,WX5817,II18008);
  nand NAND2_3123(II18007,II18009,II18010);
  nand NAND2_3124(II18015,WX5881,II18007);
  nand NAND2_3125(II18016,WX5881,II18015);
  nand NAND2_3126(II18017,II18007,II18015);
  nand NAND2_3127(II18006,II18016,II18017);
  nand NAND2_3128(II18023,WX5945,WX6009);
  nand NAND2_3129(II18024,WX5945,II18023);
  nand NAND2_3130(II18025,WX6009,II18023);
  nand NAND2_3131(II18022,II18024,II18025);
  nand NAND2_3132(II18030,II18006,II18022);
  nand NAND2_3133(II18031,II18006,II18030);
  nand NAND2_3134(II18032,II18022,II18030);
  nand NAND2_3135(WX6072,II18031,II18032);
  nand NAND2_3136(II18039,WX6173,WX5819);
  nand NAND2_3137(II18040,WX6173,II18039);
  nand NAND2_3138(II18041,WX5819,II18039);
  nand NAND2_3139(II18038,II18040,II18041);
  nand NAND2_3140(II18046,WX5883,II18038);
  nand NAND2_3141(II18047,WX5883,II18046);
  nand NAND2_3142(II18048,II18038,II18046);
  nand NAND2_3143(II18037,II18047,II18048);
  nand NAND2_3144(II18054,WX5947,WX6011);
  nand NAND2_3145(II18055,WX5947,II18054);
  nand NAND2_3146(II18056,WX6011,II18054);
  nand NAND2_3147(II18053,II18055,II18056);
  nand NAND2_3148(II18061,II18037,II18053);
  nand NAND2_3149(II18062,II18037,II18061);
  nand NAND2_3150(II18063,II18053,II18061);
  nand NAND2_3151(WX6073,II18062,II18063);
  nand NAND2_3152(II18070,WX6173,WX5821);
  nand NAND2_3153(II18071,WX6173,II18070);
  nand NAND2_3154(II18072,WX5821,II18070);
  nand NAND2_3155(II18069,II18071,II18072);
  nand NAND2_3156(II18077,WX5885,II18069);
  nand NAND2_3157(II18078,WX5885,II18077);
  nand NAND2_3158(II18079,II18069,II18077);
  nand NAND2_3159(II18068,II18078,II18079);
  nand NAND2_3160(II18085,WX5949,WX6013);
  nand NAND2_3161(II18086,WX5949,II18085);
  nand NAND2_3162(II18087,WX6013,II18085);
  nand NAND2_3163(II18084,II18086,II18087);
  nand NAND2_3164(II18092,II18068,II18084);
  nand NAND2_3165(II18093,II18068,II18092);
  nand NAND2_3166(II18094,II18084,II18092);
  nand NAND2_3167(WX6074,II18093,II18094);
  nand NAND2_3168(II18101,WX6173,WX5823);
  nand NAND2_3169(II18102,WX6173,II18101);
  nand NAND2_3170(II18103,WX5823,II18101);
  nand NAND2_3171(II18100,II18102,II18103);
  nand NAND2_3172(II18108,WX5887,II18100);
  nand NAND2_3173(II18109,WX5887,II18108);
  nand NAND2_3174(II18110,II18100,II18108);
  nand NAND2_3175(II18099,II18109,II18110);
  nand NAND2_3176(II18116,WX5951,WX6015);
  nand NAND2_3177(II18117,WX5951,II18116);
  nand NAND2_3178(II18118,WX6015,II18116);
  nand NAND2_3179(II18115,II18117,II18118);
  nand NAND2_3180(II18123,II18099,II18115);
  nand NAND2_3181(II18124,II18099,II18123);
  nand NAND2_3182(II18125,II18115,II18123);
  nand NAND2_3183(WX6075,II18124,II18125);
  nand NAND2_3184(II18132,WX6173,WX5825);
  nand NAND2_3185(II18133,WX6173,II18132);
  nand NAND2_3186(II18134,WX5825,II18132);
  nand NAND2_3187(II18131,II18133,II18134);
  nand NAND2_3188(II18139,WX5889,II18131);
  nand NAND2_3189(II18140,WX5889,II18139);
  nand NAND2_3190(II18141,II18131,II18139);
  nand NAND2_3191(II18130,II18140,II18141);
  nand NAND2_3192(II18147,WX5953,WX6017);
  nand NAND2_3193(II18148,WX5953,II18147);
  nand NAND2_3194(II18149,WX6017,II18147);
  nand NAND2_3195(II18146,II18148,II18149);
  nand NAND2_3196(II18154,II18130,II18146);
  nand NAND2_3197(II18155,II18130,II18154);
  nand NAND2_3198(II18156,II18146,II18154);
  nand NAND2_3199(WX6076,II18155,II18156);
  nand NAND2_3200(II18163,WX6173,WX5827);
  nand NAND2_3201(II18164,WX6173,II18163);
  nand NAND2_3202(II18165,WX5827,II18163);
  nand NAND2_3203(II18162,II18164,II18165);
  nand NAND2_3204(II18170,WX5891,II18162);
  nand NAND2_3205(II18171,WX5891,II18170);
  nand NAND2_3206(II18172,II18162,II18170);
  nand NAND2_3207(II18161,II18171,II18172);
  nand NAND2_3208(II18178,WX5955,WX6019);
  nand NAND2_3209(II18179,WX5955,II18178);
  nand NAND2_3210(II18180,WX6019,II18178);
  nand NAND2_3211(II18177,II18179,II18180);
  nand NAND2_3212(II18185,II18161,II18177);
  nand NAND2_3213(II18186,II18161,II18185);
  nand NAND2_3214(II18187,II18177,II18185);
  nand NAND2_3215(WX6077,II18186,II18187);
  nand NAND2_3216(II18194,WX6173,WX5829);
  nand NAND2_3217(II18195,WX6173,II18194);
  nand NAND2_3218(II18196,WX5829,II18194);
  nand NAND2_3219(II18193,II18195,II18196);
  nand NAND2_3220(II18201,WX5893,II18193);
  nand NAND2_3221(II18202,WX5893,II18201);
  nand NAND2_3222(II18203,II18193,II18201);
  nand NAND2_3223(II18192,II18202,II18203);
  nand NAND2_3224(II18209,WX5957,WX6021);
  nand NAND2_3225(II18210,WX5957,II18209);
  nand NAND2_3226(II18211,WX6021,II18209);
  nand NAND2_3227(II18208,II18210,II18211);
  nand NAND2_3228(II18216,II18192,II18208);
  nand NAND2_3229(II18217,II18192,II18216);
  nand NAND2_3230(II18218,II18208,II18216);
  nand NAND2_3231(WX6078,II18217,II18218);
  nand NAND2_3232(II18225,WX6173,WX5831);
  nand NAND2_3233(II18226,WX6173,II18225);
  nand NAND2_3234(II18227,WX5831,II18225);
  nand NAND2_3235(II18224,II18226,II18227);
  nand NAND2_3236(II18232,WX5895,II18224);
  nand NAND2_3237(II18233,WX5895,II18232);
  nand NAND2_3238(II18234,II18224,II18232);
  nand NAND2_3239(II18223,II18233,II18234);
  nand NAND2_3240(II18240,WX5959,WX6023);
  nand NAND2_3241(II18241,WX5959,II18240);
  nand NAND2_3242(II18242,WX6023,II18240);
  nand NAND2_3243(II18239,II18241,II18242);
  nand NAND2_3244(II18247,II18223,II18239);
  nand NAND2_3245(II18248,II18223,II18247);
  nand NAND2_3246(II18249,II18239,II18247);
  nand NAND2_3247(WX6079,II18248,II18249);
  nand NAND2_3248(II18256,WX6173,WX5833);
  nand NAND2_3249(II18257,WX6173,II18256);
  nand NAND2_3250(II18258,WX5833,II18256);
  nand NAND2_3251(II18255,II18257,II18258);
  nand NAND2_3252(II18263,WX5897,II18255);
  nand NAND2_3253(II18264,WX5897,II18263);
  nand NAND2_3254(II18265,II18255,II18263);
  nand NAND2_3255(II18254,II18264,II18265);
  nand NAND2_3256(II18271,WX5961,WX6025);
  nand NAND2_3257(II18272,WX5961,II18271);
  nand NAND2_3258(II18273,WX6025,II18271);
  nand NAND2_3259(II18270,II18272,II18273);
  nand NAND2_3260(II18278,II18254,II18270);
  nand NAND2_3261(II18279,II18254,II18278);
  nand NAND2_3262(II18280,II18270,II18278);
  nand NAND2_3263(WX6080,II18279,II18280);
  nand NAND2_3264(II18287,WX6173,WX5835);
  nand NAND2_3265(II18288,WX6173,II18287);
  nand NAND2_3266(II18289,WX5835,II18287);
  nand NAND2_3267(II18286,II18288,II18289);
  nand NAND2_3268(II18294,WX5899,II18286);
  nand NAND2_3269(II18295,WX5899,II18294);
  nand NAND2_3270(II18296,II18286,II18294);
  nand NAND2_3271(II18285,II18295,II18296);
  nand NAND2_3272(II18302,WX5963,WX6027);
  nand NAND2_3273(II18303,WX5963,II18302);
  nand NAND2_3274(II18304,WX6027,II18302);
  nand NAND2_3275(II18301,II18303,II18304);
  nand NAND2_3276(II18309,II18285,II18301);
  nand NAND2_3277(II18310,II18285,II18309);
  nand NAND2_3278(II18311,II18301,II18309);
  nand NAND2_3279(WX6081,II18310,II18311);
  nand NAND2_3280(II18318,WX6173,WX5837);
  nand NAND2_3281(II18319,WX6173,II18318);
  nand NAND2_3282(II18320,WX5837,II18318);
  nand NAND2_3283(II18317,II18319,II18320);
  nand NAND2_3284(II18325,WX5901,II18317);
  nand NAND2_3285(II18326,WX5901,II18325);
  nand NAND2_3286(II18327,II18317,II18325);
  nand NAND2_3287(II18316,II18326,II18327);
  nand NAND2_3288(II18333,WX5965,WX6029);
  nand NAND2_3289(II18334,WX5965,II18333);
  nand NAND2_3290(II18335,WX6029,II18333);
  nand NAND2_3291(II18332,II18334,II18335);
  nand NAND2_3292(II18340,II18316,II18332);
  nand NAND2_3293(II18341,II18316,II18340);
  nand NAND2_3294(II18342,II18332,II18340);
  nand NAND2_3295(WX6082,II18341,II18342);
  nand NAND2_3296(II18349,WX6173,WX5839);
  nand NAND2_3297(II18350,WX6173,II18349);
  nand NAND2_3298(II18351,WX5839,II18349);
  nand NAND2_3299(II18348,II18350,II18351);
  nand NAND2_3300(II18356,WX5903,II18348);
  nand NAND2_3301(II18357,WX5903,II18356);
  nand NAND2_3302(II18358,II18348,II18356);
  nand NAND2_3303(II18347,II18357,II18358);
  nand NAND2_3304(II18364,WX5967,WX6031);
  nand NAND2_3305(II18365,WX5967,II18364);
  nand NAND2_3306(II18366,WX6031,II18364);
  nand NAND2_3307(II18363,II18365,II18366);
  nand NAND2_3308(II18371,II18347,II18363);
  nand NAND2_3309(II18372,II18347,II18371);
  nand NAND2_3310(II18373,II18363,II18371);
  nand NAND2_3311(WX6083,II18372,II18373);
  nand NAND2_3312(II18380,WX6173,WX5841);
  nand NAND2_3313(II18381,WX6173,II18380);
  nand NAND2_3314(II18382,WX5841,II18380);
  nand NAND2_3315(II18379,II18381,II18382);
  nand NAND2_3316(II18387,WX5905,II18379);
  nand NAND2_3317(II18388,WX5905,II18387);
  nand NAND2_3318(II18389,II18379,II18387);
  nand NAND2_3319(II18378,II18388,II18389);
  nand NAND2_3320(II18395,WX5969,WX6033);
  nand NAND2_3321(II18396,WX5969,II18395);
  nand NAND2_3322(II18397,WX6033,II18395);
  nand NAND2_3323(II18394,II18396,II18397);
  nand NAND2_3324(II18402,II18378,II18394);
  nand NAND2_3325(II18403,II18378,II18402);
  nand NAND2_3326(II18404,II18394,II18402);
  nand NAND2_3327(WX6084,II18403,II18404);
  nand NAND2_3328(II18411,WX6173,WX5843);
  nand NAND2_3329(II18412,WX6173,II18411);
  nand NAND2_3330(II18413,WX5843,II18411);
  nand NAND2_3331(II18410,II18412,II18413);
  nand NAND2_3332(II18418,WX5907,II18410);
  nand NAND2_3333(II18419,WX5907,II18418);
  nand NAND2_3334(II18420,II18410,II18418);
  nand NAND2_3335(II18409,II18419,II18420);
  nand NAND2_3336(II18426,WX5971,WX6035);
  nand NAND2_3337(II18427,WX5971,II18426);
  nand NAND2_3338(II18428,WX6035,II18426);
  nand NAND2_3339(II18425,II18427,II18428);
  nand NAND2_3340(II18433,II18409,II18425);
  nand NAND2_3341(II18434,II18409,II18433);
  nand NAND2_3342(II18435,II18425,II18433);
  nand NAND2_3343(WX6085,II18434,II18435);
  nand NAND2_3344(II18442,WX6173,WX5845);
  nand NAND2_3345(II18443,WX6173,II18442);
  nand NAND2_3346(II18444,WX5845,II18442);
  nand NAND2_3347(II18441,II18443,II18444);
  nand NAND2_3348(II18449,WX5909,II18441);
  nand NAND2_3349(II18450,WX5909,II18449);
  nand NAND2_3350(II18451,II18441,II18449);
  nand NAND2_3351(II18440,II18450,II18451);
  nand NAND2_3352(II18457,WX5973,WX6037);
  nand NAND2_3353(II18458,WX5973,II18457);
  nand NAND2_3354(II18459,WX6037,II18457);
  nand NAND2_3355(II18456,II18458,II18459);
  nand NAND2_3356(II18464,II18440,II18456);
  nand NAND2_3357(II18465,II18440,II18464);
  nand NAND2_3358(II18466,II18456,II18464);
  nand NAND2_3359(WX6086,II18465,II18466);
  nand NAND2_3360(II18473,WX6173,WX5847);
  nand NAND2_3361(II18474,WX6173,II18473);
  nand NAND2_3362(II18475,WX5847,II18473);
  nand NAND2_3363(II18472,II18474,II18475);
  nand NAND2_3364(II18480,WX5911,II18472);
  nand NAND2_3365(II18481,WX5911,II18480);
  nand NAND2_3366(II18482,II18472,II18480);
  nand NAND2_3367(II18471,II18481,II18482);
  nand NAND2_3368(II18488,WX5975,WX6039);
  nand NAND2_3369(II18489,WX5975,II18488);
  nand NAND2_3370(II18490,WX6039,II18488);
  nand NAND2_3371(II18487,II18489,II18490);
  nand NAND2_3372(II18495,II18471,II18487);
  nand NAND2_3373(II18496,II18471,II18495);
  nand NAND2_3374(II18497,II18487,II18495);
  nand NAND2_3375(WX6087,II18496,II18497);
  nand NAND2_3376(II18504,WX6174,WX5849);
  nand NAND2_3377(II18505,WX6174,II18504);
  nand NAND2_3378(II18506,WX5849,II18504);
  nand NAND2_3379(II18503,II18505,II18506);
  nand NAND2_3380(II18511,WX5913,II18503);
  nand NAND2_3381(II18512,WX5913,II18511);
  nand NAND2_3382(II18513,II18503,II18511);
  nand NAND2_3383(II18502,II18512,II18513);
  nand NAND2_3384(II18519,WX5977,WX6041);
  nand NAND2_3385(II18520,WX5977,II18519);
  nand NAND2_3386(II18521,WX6041,II18519);
  nand NAND2_3387(II18518,II18520,II18521);
  nand NAND2_3388(II18526,II18502,II18518);
  nand NAND2_3389(II18527,II18502,II18526);
  nand NAND2_3390(II18528,II18518,II18526);
  nand NAND2_3391(WX6088,II18527,II18528);
  nand NAND2_3392(II18535,WX6174,WX5851);
  nand NAND2_3393(II18536,WX6174,II18535);
  nand NAND2_3394(II18537,WX5851,II18535);
  nand NAND2_3395(II18534,II18536,II18537);
  nand NAND2_3396(II18542,WX5915,II18534);
  nand NAND2_3397(II18543,WX5915,II18542);
  nand NAND2_3398(II18544,II18534,II18542);
  nand NAND2_3399(II18533,II18543,II18544);
  nand NAND2_3400(II18550,WX5979,WX6043);
  nand NAND2_3401(II18551,WX5979,II18550);
  nand NAND2_3402(II18552,WX6043,II18550);
  nand NAND2_3403(II18549,II18551,II18552);
  nand NAND2_3404(II18557,II18533,II18549);
  nand NAND2_3405(II18558,II18533,II18557);
  nand NAND2_3406(II18559,II18549,II18557);
  nand NAND2_3407(WX6089,II18558,II18559);
  nand NAND2_3408(II18566,WX6174,WX5853);
  nand NAND2_3409(II18567,WX6174,II18566);
  nand NAND2_3410(II18568,WX5853,II18566);
  nand NAND2_3411(II18565,II18567,II18568);
  nand NAND2_3412(II18573,WX5917,II18565);
  nand NAND2_3413(II18574,WX5917,II18573);
  nand NAND2_3414(II18575,II18565,II18573);
  nand NAND2_3415(II18564,II18574,II18575);
  nand NAND2_3416(II18581,WX5981,WX6045);
  nand NAND2_3417(II18582,WX5981,II18581);
  nand NAND2_3418(II18583,WX6045,II18581);
  nand NAND2_3419(II18580,II18582,II18583);
  nand NAND2_3420(II18588,II18564,II18580);
  nand NAND2_3421(II18589,II18564,II18588);
  nand NAND2_3422(II18590,II18580,II18588);
  nand NAND2_3423(WX6090,II18589,II18590);
  nand NAND2_3424(II18597,WX6174,WX5855);
  nand NAND2_3425(II18598,WX6174,II18597);
  nand NAND2_3426(II18599,WX5855,II18597);
  nand NAND2_3427(II18596,II18598,II18599);
  nand NAND2_3428(II18604,WX5919,II18596);
  nand NAND2_3429(II18605,WX5919,II18604);
  nand NAND2_3430(II18606,II18596,II18604);
  nand NAND2_3431(II18595,II18605,II18606);
  nand NAND2_3432(II18612,WX5983,WX6047);
  nand NAND2_3433(II18613,WX5983,II18612);
  nand NAND2_3434(II18614,WX6047,II18612);
  nand NAND2_3435(II18611,II18613,II18614);
  nand NAND2_3436(II18619,II18595,II18611);
  nand NAND2_3437(II18620,II18595,II18619);
  nand NAND2_3438(II18621,II18611,II18619);
  nand NAND2_3439(WX6091,II18620,II18621);
  nand NAND2_3440(II18628,WX6174,WX5857);
  nand NAND2_3441(II18629,WX6174,II18628);
  nand NAND2_3442(II18630,WX5857,II18628);
  nand NAND2_3443(II18627,II18629,II18630);
  nand NAND2_3444(II18635,WX5921,II18627);
  nand NAND2_3445(II18636,WX5921,II18635);
  nand NAND2_3446(II18637,II18627,II18635);
  nand NAND2_3447(II18626,II18636,II18637);
  nand NAND2_3448(II18643,WX5985,WX6049);
  nand NAND2_3449(II18644,WX5985,II18643);
  nand NAND2_3450(II18645,WX6049,II18643);
  nand NAND2_3451(II18642,II18644,II18645);
  nand NAND2_3452(II18650,II18626,II18642);
  nand NAND2_3453(II18651,II18626,II18650);
  nand NAND2_3454(II18652,II18642,II18650);
  nand NAND2_3455(WX6092,II18651,II18652);
  nand NAND2_3456(II18659,WX6174,WX5859);
  nand NAND2_3457(II18660,WX6174,II18659);
  nand NAND2_3458(II18661,WX5859,II18659);
  nand NAND2_3459(II18658,II18660,II18661);
  nand NAND2_3460(II18666,WX5923,II18658);
  nand NAND2_3461(II18667,WX5923,II18666);
  nand NAND2_3462(II18668,II18658,II18666);
  nand NAND2_3463(II18657,II18667,II18668);
  nand NAND2_3464(II18674,WX5987,WX6051);
  nand NAND2_3465(II18675,WX5987,II18674);
  nand NAND2_3466(II18676,WX6051,II18674);
  nand NAND2_3467(II18673,II18675,II18676);
  nand NAND2_3468(II18681,II18657,II18673);
  nand NAND2_3469(II18682,II18657,II18681);
  nand NAND2_3470(II18683,II18673,II18681);
  nand NAND2_3471(WX6093,II18682,II18683);
  nand NAND2_3472(II18690,WX6174,WX5861);
  nand NAND2_3473(II18691,WX6174,II18690);
  nand NAND2_3474(II18692,WX5861,II18690);
  nand NAND2_3475(II18689,II18691,II18692);
  nand NAND2_3476(II18697,WX5925,II18689);
  nand NAND2_3477(II18698,WX5925,II18697);
  nand NAND2_3478(II18699,II18689,II18697);
  nand NAND2_3479(II18688,II18698,II18699);
  nand NAND2_3480(II18705,WX5989,WX6053);
  nand NAND2_3481(II18706,WX5989,II18705);
  nand NAND2_3482(II18707,WX6053,II18705);
  nand NAND2_3483(II18704,II18706,II18707);
  nand NAND2_3484(II18712,II18688,II18704);
  nand NAND2_3485(II18713,II18688,II18712);
  nand NAND2_3486(II18714,II18704,II18712);
  nand NAND2_3487(WX6094,II18713,II18714);
  nand NAND2_3488(II18721,WX6174,WX5863);
  nand NAND2_3489(II18722,WX6174,II18721);
  nand NAND2_3490(II18723,WX5863,II18721);
  nand NAND2_3491(II18720,II18722,II18723);
  nand NAND2_3492(II18728,WX5927,II18720);
  nand NAND2_3493(II18729,WX5927,II18728);
  nand NAND2_3494(II18730,II18720,II18728);
  nand NAND2_3495(II18719,II18729,II18730);
  nand NAND2_3496(II18736,WX5991,WX6055);
  nand NAND2_3497(II18737,WX5991,II18736);
  nand NAND2_3498(II18738,WX6055,II18736);
  nand NAND2_3499(II18735,II18737,II18738);
  nand NAND2_3500(II18743,II18719,II18735);
  nand NAND2_3501(II18744,II18719,II18743);
  nand NAND2_3502(II18745,II18735,II18743);
  nand NAND2_3503(WX6095,II18744,II18745);
  nand NAND2_3504(II18752,WX6174,WX5865);
  nand NAND2_3505(II18753,WX6174,II18752);
  nand NAND2_3506(II18754,WX5865,II18752);
  nand NAND2_3507(II18751,II18753,II18754);
  nand NAND2_3508(II18759,WX5929,II18751);
  nand NAND2_3509(II18760,WX5929,II18759);
  nand NAND2_3510(II18761,II18751,II18759);
  nand NAND2_3511(II18750,II18760,II18761);
  nand NAND2_3512(II18767,WX5993,WX6057);
  nand NAND2_3513(II18768,WX5993,II18767);
  nand NAND2_3514(II18769,WX6057,II18767);
  nand NAND2_3515(II18766,II18768,II18769);
  nand NAND2_3516(II18774,II18750,II18766);
  nand NAND2_3517(II18775,II18750,II18774);
  nand NAND2_3518(II18776,II18766,II18774);
  nand NAND2_3519(WX6096,II18775,II18776);
  nand NAND2_3520(II18783,WX6174,WX5867);
  nand NAND2_3521(II18784,WX6174,II18783);
  nand NAND2_3522(II18785,WX5867,II18783);
  nand NAND2_3523(II18782,II18784,II18785);
  nand NAND2_3524(II18790,WX5931,II18782);
  nand NAND2_3525(II18791,WX5931,II18790);
  nand NAND2_3526(II18792,II18782,II18790);
  nand NAND2_3527(II18781,II18791,II18792);
  nand NAND2_3528(II18798,WX5995,WX6059);
  nand NAND2_3529(II18799,WX5995,II18798);
  nand NAND2_3530(II18800,WX6059,II18798);
  nand NAND2_3531(II18797,II18799,II18800);
  nand NAND2_3532(II18805,II18781,II18797);
  nand NAND2_3533(II18806,II18781,II18805);
  nand NAND2_3534(II18807,II18797,II18805);
  nand NAND2_3535(WX6097,II18806,II18807);
  nand NAND2_3536(II18814,WX6174,WX5869);
  nand NAND2_3537(II18815,WX6174,II18814);
  nand NAND2_3538(II18816,WX5869,II18814);
  nand NAND2_3539(II18813,II18815,II18816);
  nand NAND2_3540(II18821,WX5933,II18813);
  nand NAND2_3541(II18822,WX5933,II18821);
  nand NAND2_3542(II18823,II18813,II18821);
  nand NAND2_3543(II18812,II18822,II18823);
  nand NAND2_3544(II18829,WX5997,WX6061);
  nand NAND2_3545(II18830,WX5997,II18829);
  nand NAND2_3546(II18831,WX6061,II18829);
  nand NAND2_3547(II18828,II18830,II18831);
  nand NAND2_3548(II18836,II18812,II18828);
  nand NAND2_3549(II18837,II18812,II18836);
  nand NAND2_3550(II18838,II18828,II18836);
  nand NAND2_3551(WX6098,II18837,II18838);
  nand NAND2_3552(II18845,WX6174,WX5871);
  nand NAND2_3553(II18846,WX6174,II18845);
  nand NAND2_3554(II18847,WX5871,II18845);
  nand NAND2_3555(II18844,II18846,II18847);
  nand NAND2_3556(II18852,WX5935,II18844);
  nand NAND2_3557(II18853,WX5935,II18852);
  nand NAND2_3558(II18854,II18844,II18852);
  nand NAND2_3559(II18843,II18853,II18854);
  nand NAND2_3560(II18860,WX5999,WX6063);
  nand NAND2_3561(II18861,WX5999,II18860);
  nand NAND2_3562(II18862,WX6063,II18860);
  nand NAND2_3563(II18859,II18861,II18862);
  nand NAND2_3564(II18867,II18843,II18859);
  nand NAND2_3565(II18868,II18843,II18867);
  nand NAND2_3566(II18869,II18859,II18867);
  nand NAND2_3567(WX6099,II18868,II18869);
  nand NAND2_3568(II18876,WX6174,WX5873);
  nand NAND2_3569(II18877,WX6174,II18876);
  nand NAND2_3570(II18878,WX5873,II18876);
  nand NAND2_3571(II18875,II18877,II18878);
  nand NAND2_3572(II18883,WX5937,II18875);
  nand NAND2_3573(II18884,WX5937,II18883);
  nand NAND2_3574(II18885,II18875,II18883);
  nand NAND2_3575(II18874,II18884,II18885);
  nand NAND2_3576(II18891,WX6001,WX6065);
  nand NAND2_3577(II18892,WX6001,II18891);
  nand NAND2_3578(II18893,WX6065,II18891);
  nand NAND2_3579(II18890,II18892,II18893);
  nand NAND2_3580(II18898,II18874,II18890);
  nand NAND2_3581(II18899,II18874,II18898);
  nand NAND2_3582(II18900,II18890,II18898);
  nand NAND2_3583(WX6100,II18899,II18900);
  nand NAND2_3584(II18907,WX6174,WX5875);
  nand NAND2_3585(II18908,WX6174,II18907);
  nand NAND2_3586(II18909,WX5875,II18907);
  nand NAND2_3587(II18906,II18908,II18909);
  nand NAND2_3588(II18914,WX5939,II18906);
  nand NAND2_3589(II18915,WX5939,II18914);
  nand NAND2_3590(II18916,II18906,II18914);
  nand NAND2_3591(II18905,II18915,II18916);
  nand NAND2_3592(II18922,WX6003,WX6067);
  nand NAND2_3593(II18923,WX6003,II18922);
  nand NAND2_3594(II18924,WX6067,II18922);
  nand NAND2_3595(II18921,II18923,II18924);
  nand NAND2_3596(II18929,II18905,II18921);
  nand NAND2_3597(II18930,II18905,II18929);
  nand NAND2_3598(II18931,II18921,II18929);
  nand NAND2_3599(WX6101,II18930,II18931);
  nand NAND2_3600(II18938,WX6174,WX5877);
  nand NAND2_3601(II18939,WX6174,II18938);
  nand NAND2_3602(II18940,WX5877,II18938);
  nand NAND2_3603(II18937,II18939,II18940);
  nand NAND2_3604(II18945,WX5941,II18937);
  nand NAND2_3605(II18946,WX5941,II18945);
  nand NAND2_3606(II18947,II18937,II18945);
  nand NAND2_3607(II18936,II18946,II18947);
  nand NAND2_3608(II18953,WX6005,WX6069);
  nand NAND2_3609(II18954,WX6005,II18953);
  nand NAND2_3610(II18955,WX6069,II18953);
  nand NAND2_3611(II18952,II18954,II18955);
  nand NAND2_3612(II18960,II18936,II18952);
  nand NAND2_3613(II18961,II18936,II18960);
  nand NAND2_3614(II18962,II18952,II18960);
  nand NAND2_3615(WX6102,II18961,II18962);
  nand NAND2_3616(II18969,WX6174,WX5879);
  nand NAND2_3617(II18970,WX6174,II18969);
  nand NAND2_3618(II18971,WX5879,II18969);
  nand NAND2_3619(II18968,II18970,II18971);
  nand NAND2_3620(II18976,WX5943,II18968);
  nand NAND2_3621(II18977,WX5943,II18976);
  nand NAND2_3622(II18978,II18968,II18976);
  nand NAND2_3623(II18967,II18977,II18978);
  nand NAND2_3624(II18984,WX6007,WX6071);
  nand NAND2_3625(II18985,WX6007,II18984);
  nand NAND2_3626(II18986,WX6071,II18984);
  nand NAND2_3627(II18983,II18985,II18986);
  nand NAND2_3628(II18991,II18967,II18983);
  nand NAND2_3629(II18992,II18967,II18991);
  nand NAND2_3630(II18993,II18983,II18991);
  nand NAND2_3631(WX6103,II18992,II18993);
  nand NAND2_3632(II19072,WX5752,WX5657);
  nand NAND2_3633(II19073,WX5752,II19072);
  nand NAND2_3634(II19074,WX5657,II19072);
  nand NAND2_3635(WX6178,II19073,II19074);
  nand NAND2_3636(II19085,WX5753,WX5659);
  nand NAND2_3637(II19086,WX5753,II19085);
  nand NAND2_3638(II19087,WX5659,II19085);
  nand NAND2_3639(WX6185,II19086,II19087);
  nand NAND2_3640(II19098,WX5754,WX5661);
  nand NAND2_3641(II19099,WX5754,II19098);
  nand NAND2_3642(II19100,WX5661,II19098);
  nand NAND2_3643(WX6192,II19099,II19100);
  nand NAND2_3644(II19111,WX5755,WX5663);
  nand NAND2_3645(II19112,WX5755,II19111);
  nand NAND2_3646(II19113,WX5663,II19111);
  nand NAND2_3647(WX6199,II19112,II19113);
  nand NAND2_3648(II19124,WX5756,WX5665);
  nand NAND2_3649(II19125,WX5756,II19124);
  nand NAND2_3650(II19126,WX5665,II19124);
  nand NAND2_3651(WX6206,II19125,II19126);
  nand NAND2_3652(II19137,WX5757,WX5667);
  nand NAND2_3653(II19138,WX5757,II19137);
  nand NAND2_3654(II19139,WX5667,II19137);
  nand NAND2_3655(WX6213,II19138,II19139);
  nand NAND2_3656(II19150,WX5758,WX5669);
  nand NAND2_3657(II19151,WX5758,II19150);
  nand NAND2_3658(II19152,WX5669,II19150);
  nand NAND2_3659(WX6220,II19151,II19152);
  nand NAND2_3660(II19163,WX5759,WX5671);
  nand NAND2_3661(II19164,WX5759,II19163);
  nand NAND2_3662(II19165,WX5671,II19163);
  nand NAND2_3663(WX6227,II19164,II19165);
  nand NAND2_3664(II19176,WX5760,WX5673);
  nand NAND2_3665(II19177,WX5760,II19176);
  nand NAND2_3666(II19178,WX5673,II19176);
  nand NAND2_3667(WX6234,II19177,II19178);
  nand NAND2_3668(II19189,WX5761,WX5675);
  nand NAND2_3669(II19190,WX5761,II19189);
  nand NAND2_3670(II19191,WX5675,II19189);
  nand NAND2_3671(WX6241,II19190,II19191);
  nand NAND2_3672(II19202,WX5762,WX5677);
  nand NAND2_3673(II19203,WX5762,II19202);
  nand NAND2_3674(II19204,WX5677,II19202);
  nand NAND2_3675(WX6248,II19203,II19204);
  nand NAND2_3676(II19215,WX5763,WX5679);
  nand NAND2_3677(II19216,WX5763,II19215);
  nand NAND2_3678(II19217,WX5679,II19215);
  nand NAND2_3679(WX6255,II19216,II19217);
  nand NAND2_3680(II19228,WX5764,WX5681);
  nand NAND2_3681(II19229,WX5764,II19228);
  nand NAND2_3682(II19230,WX5681,II19228);
  nand NAND2_3683(WX6262,II19229,II19230);
  nand NAND2_3684(II19241,WX5765,WX5683);
  nand NAND2_3685(II19242,WX5765,II19241);
  nand NAND2_3686(II19243,WX5683,II19241);
  nand NAND2_3687(WX6269,II19242,II19243);
  nand NAND2_3688(II19254,WX5766,WX5685);
  nand NAND2_3689(II19255,WX5766,II19254);
  nand NAND2_3690(II19256,WX5685,II19254);
  nand NAND2_3691(WX6276,II19255,II19256);
  nand NAND2_3692(II19267,WX5767,WX5687);
  nand NAND2_3693(II19268,WX5767,II19267);
  nand NAND2_3694(II19269,WX5687,II19267);
  nand NAND2_3695(WX6283,II19268,II19269);
  nand NAND2_3696(II19280,WX5768,WX5689);
  nand NAND2_3697(II19281,WX5768,II19280);
  nand NAND2_3698(II19282,WX5689,II19280);
  nand NAND2_3699(WX6290,II19281,II19282);
  nand NAND2_3700(II19293,WX5769,WX5691);
  nand NAND2_3701(II19294,WX5769,II19293);
  nand NAND2_3702(II19295,WX5691,II19293);
  nand NAND2_3703(WX6297,II19294,II19295);
  nand NAND2_3704(II19306,WX5770,WX5693);
  nand NAND2_3705(II19307,WX5770,II19306);
  nand NAND2_3706(II19308,WX5693,II19306);
  nand NAND2_3707(WX6304,II19307,II19308);
  nand NAND2_3708(II19319,WX5771,WX5695);
  nand NAND2_3709(II19320,WX5771,II19319);
  nand NAND2_3710(II19321,WX5695,II19319);
  nand NAND2_3711(WX6311,II19320,II19321);
  nand NAND2_3712(II19332,WX5772,WX5697);
  nand NAND2_3713(II19333,WX5772,II19332);
  nand NAND2_3714(II19334,WX5697,II19332);
  nand NAND2_3715(WX6318,II19333,II19334);
  nand NAND2_3716(II19345,WX5773,WX5699);
  nand NAND2_3717(II19346,WX5773,II19345);
  nand NAND2_3718(II19347,WX5699,II19345);
  nand NAND2_3719(WX6325,II19346,II19347);
  nand NAND2_3720(II19358,WX5774,WX5701);
  nand NAND2_3721(II19359,WX5774,II19358);
  nand NAND2_3722(II19360,WX5701,II19358);
  nand NAND2_3723(WX6332,II19359,II19360);
  nand NAND2_3724(II19371,WX5775,WX5703);
  nand NAND2_3725(II19372,WX5775,II19371);
  nand NAND2_3726(II19373,WX5703,II19371);
  nand NAND2_3727(WX6339,II19372,II19373);
  nand NAND2_3728(II19384,WX5776,WX5705);
  nand NAND2_3729(II19385,WX5776,II19384);
  nand NAND2_3730(II19386,WX5705,II19384);
  nand NAND2_3731(WX6346,II19385,II19386);
  nand NAND2_3732(II19397,WX5777,WX5707);
  nand NAND2_3733(II19398,WX5777,II19397);
  nand NAND2_3734(II19399,WX5707,II19397);
  nand NAND2_3735(WX6353,II19398,II19399);
  nand NAND2_3736(II19410,WX5778,WX5709);
  nand NAND2_3737(II19411,WX5778,II19410);
  nand NAND2_3738(II19412,WX5709,II19410);
  nand NAND2_3739(WX6360,II19411,II19412);
  nand NAND2_3740(II19423,WX5779,WX5711);
  nand NAND2_3741(II19424,WX5779,II19423);
  nand NAND2_3742(II19425,WX5711,II19423);
  nand NAND2_3743(WX6367,II19424,II19425);
  nand NAND2_3744(II19436,WX5780,WX5713);
  nand NAND2_3745(II19437,WX5780,II19436);
  nand NAND2_3746(II19438,WX5713,II19436);
  nand NAND2_3747(WX6374,II19437,II19438);
  nand NAND2_3748(II19449,WX5781,WX5715);
  nand NAND2_3749(II19450,WX5781,II19449);
  nand NAND2_3750(II19451,WX5715,II19449);
  nand NAND2_3751(WX6381,II19450,II19451);
  nand NAND2_3752(II19462,WX5782,WX5717);
  nand NAND2_3753(II19463,WX5782,II19462);
  nand NAND2_3754(II19464,WX5717,II19462);
  nand NAND2_3755(WX6388,II19463,II19464);
  nand NAND2_3756(II19475,WX5783,WX5719);
  nand NAND2_3757(II19476,WX5783,II19475);
  nand NAND2_3758(II19477,WX5719,II19475);
  nand NAND2_3759(WX6395,II19476,II19477);
  nand NAND2_3760(II19490,WX5799,CRC_OUT_5_31);
  nand NAND2_3761(II19491,WX5799,II19490);
  nand NAND2_3762(II19492,CRC_OUT_5_31,II19490);
  nand NAND2_3763(II19489,II19491,II19492);
  nand NAND2_3764(II19497,CRC_OUT_5_15,II19489);
  nand NAND2_3765(II19498,CRC_OUT_5_15,II19497);
  nand NAND2_3766(II19499,II19489,II19497);
  nand NAND2_3767(WX6403,II19498,II19499);
  nand NAND2_3768(II19505,WX5804,CRC_OUT_5_31);
  nand NAND2_3769(II19506,WX5804,II19505);
  nand NAND2_3770(II19507,CRC_OUT_5_31,II19505);
  nand NAND2_3771(II19504,II19506,II19507);
  nand NAND2_3772(II19512,CRC_OUT_5_10,II19504);
  nand NAND2_3773(II19513,CRC_OUT_5_10,II19512);
  nand NAND2_3774(II19514,II19504,II19512);
  nand NAND2_3775(WX6404,II19513,II19514);
  nand NAND2_3776(II19520,WX5811,CRC_OUT_5_31);
  nand NAND2_3777(II19521,WX5811,II19520);
  nand NAND2_3778(II19522,CRC_OUT_5_31,II19520);
  nand NAND2_3779(II19519,II19521,II19522);
  nand NAND2_3780(II19527,CRC_OUT_5_3,II19519);
  nand NAND2_3781(II19528,CRC_OUT_5_3,II19527);
  nand NAND2_3782(II19529,II19519,II19527);
  nand NAND2_3783(WX6405,II19528,II19529);
  nand NAND2_3784(II19534,WX5815,CRC_OUT_5_31);
  nand NAND2_3785(II19535,WX5815,II19534);
  nand NAND2_3786(II19536,CRC_OUT_5_31,II19534);
  nand NAND2_3787(WX6406,II19535,II19536);
  nand NAND2_3788(II19541,WX5784,CRC_OUT_5_30);
  nand NAND2_3789(II19542,WX5784,II19541);
  nand NAND2_3790(II19543,CRC_OUT_5_30,II19541);
  nand NAND2_3791(WX6407,II19542,II19543);
  nand NAND2_3792(II19548,WX5785,CRC_OUT_5_29);
  nand NAND2_3793(II19549,WX5785,II19548);
  nand NAND2_3794(II19550,CRC_OUT_5_29,II19548);
  nand NAND2_3795(WX6408,II19549,II19550);
  nand NAND2_3796(II19555,WX5786,CRC_OUT_5_28);
  nand NAND2_3797(II19556,WX5786,II19555);
  nand NAND2_3798(II19557,CRC_OUT_5_28,II19555);
  nand NAND2_3799(WX6409,II19556,II19557);
  nand NAND2_3800(II19562,WX5787,CRC_OUT_5_27);
  nand NAND2_3801(II19563,WX5787,II19562);
  nand NAND2_3802(II19564,CRC_OUT_5_27,II19562);
  nand NAND2_3803(WX6410,II19563,II19564);
  nand NAND2_3804(II19569,WX5788,CRC_OUT_5_26);
  nand NAND2_3805(II19570,WX5788,II19569);
  nand NAND2_3806(II19571,CRC_OUT_5_26,II19569);
  nand NAND2_3807(WX6411,II19570,II19571);
  nand NAND2_3808(II19576,WX5789,CRC_OUT_5_25);
  nand NAND2_3809(II19577,WX5789,II19576);
  nand NAND2_3810(II19578,CRC_OUT_5_25,II19576);
  nand NAND2_3811(WX6412,II19577,II19578);
  nand NAND2_3812(II19583,WX5790,CRC_OUT_5_24);
  nand NAND2_3813(II19584,WX5790,II19583);
  nand NAND2_3814(II19585,CRC_OUT_5_24,II19583);
  nand NAND2_3815(WX6413,II19584,II19585);
  nand NAND2_3816(II19590,WX5791,CRC_OUT_5_23);
  nand NAND2_3817(II19591,WX5791,II19590);
  nand NAND2_3818(II19592,CRC_OUT_5_23,II19590);
  nand NAND2_3819(WX6414,II19591,II19592);
  nand NAND2_3820(II19597,WX5792,CRC_OUT_5_22);
  nand NAND2_3821(II19598,WX5792,II19597);
  nand NAND2_3822(II19599,CRC_OUT_5_22,II19597);
  nand NAND2_3823(WX6415,II19598,II19599);
  nand NAND2_3824(II19604,WX5793,CRC_OUT_5_21);
  nand NAND2_3825(II19605,WX5793,II19604);
  nand NAND2_3826(II19606,CRC_OUT_5_21,II19604);
  nand NAND2_3827(WX6416,II19605,II19606);
  nand NAND2_3828(II19611,WX5794,CRC_OUT_5_20);
  nand NAND2_3829(II19612,WX5794,II19611);
  nand NAND2_3830(II19613,CRC_OUT_5_20,II19611);
  nand NAND2_3831(WX6417,II19612,II19613);
  nand NAND2_3832(II19618,WX5795,CRC_OUT_5_19);
  nand NAND2_3833(II19619,WX5795,II19618);
  nand NAND2_3834(II19620,CRC_OUT_5_19,II19618);
  nand NAND2_3835(WX6418,II19619,II19620);
  nand NAND2_3836(II19625,WX5796,CRC_OUT_5_18);
  nand NAND2_3837(II19626,WX5796,II19625);
  nand NAND2_3838(II19627,CRC_OUT_5_18,II19625);
  nand NAND2_3839(WX6419,II19626,II19627);
  nand NAND2_3840(II19632,WX5797,CRC_OUT_5_17);
  nand NAND2_3841(II19633,WX5797,II19632);
  nand NAND2_3842(II19634,CRC_OUT_5_17,II19632);
  nand NAND2_3843(WX6420,II19633,II19634);
  nand NAND2_3844(II19639,WX5798,CRC_OUT_5_16);
  nand NAND2_3845(II19640,WX5798,II19639);
  nand NAND2_3846(II19641,CRC_OUT_5_16,II19639);
  nand NAND2_3847(WX6421,II19640,II19641);
  nand NAND2_3848(II19646,WX5800,CRC_OUT_5_14);
  nand NAND2_3849(II19647,WX5800,II19646);
  nand NAND2_3850(II19648,CRC_OUT_5_14,II19646);
  nand NAND2_3851(WX6422,II19647,II19648);
  nand NAND2_3852(II19653,WX5801,CRC_OUT_5_13);
  nand NAND2_3853(II19654,WX5801,II19653);
  nand NAND2_3854(II19655,CRC_OUT_5_13,II19653);
  nand NAND2_3855(WX6423,II19654,II19655);
  nand NAND2_3856(II19660,WX5802,CRC_OUT_5_12);
  nand NAND2_3857(II19661,WX5802,II19660);
  nand NAND2_3858(II19662,CRC_OUT_5_12,II19660);
  nand NAND2_3859(WX6424,II19661,II19662);
  nand NAND2_3860(II19667,WX5803,CRC_OUT_5_11);
  nand NAND2_3861(II19668,WX5803,II19667);
  nand NAND2_3862(II19669,CRC_OUT_5_11,II19667);
  nand NAND2_3863(WX6425,II19668,II19669);
  nand NAND2_3864(II19674,WX5805,CRC_OUT_5_9);
  nand NAND2_3865(II19675,WX5805,II19674);
  nand NAND2_3866(II19676,CRC_OUT_5_9,II19674);
  nand NAND2_3867(WX6426,II19675,II19676);
  nand NAND2_3868(II19681,WX5806,CRC_OUT_5_8);
  nand NAND2_3869(II19682,WX5806,II19681);
  nand NAND2_3870(II19683,CRC_OUT_5_8,II19681);
  nand NAND2_3871(WX6427,II19682,II19683);
  nand NAND2_3872(II19688,WX5807,CRC_OUT_5_7);
  nand NAND2_3873(II19689,WX5807,II19688);
  nand NAND2_3874(II19690,CRC_OUT_5_7,II19688);
  nand NAND2_3875(WX6428,II19689,II19690);
  nand NAND2_3876(II19695,WX5808,CRC_OUT_5_6);
  nand NAND2_3877(II19696,WX5808,II19695);
  nand NAND2_3878(II19697,CRC_OUT_5_6,II19695);
  nand NAND2_3879(WX6429,II19696,II19697);
  nand NAND2_3880(II19702,WX5809,CRC_OUT_5_5);
  nand NAND2_3881(II19703,WX5809,II19702);
  nand NAND2_3882(II19704,CRC_OUT_5_5,II19702);
  nand NAND2_3883(WX6430,II19703,II19704);
  nand NAND2_3884(II19709,WX5810,CRC_OUT_5_4);
  nand NAND2_3885(II19710,WX5810,II19709);
  nand NAND2_3886(II19711,CRC_OUT_5_4,II19709);
  nand NAND2_3887(WX6431,II19710,II19711);
  nand NAND2_3888(II19716,WX5812,CRC_OUT_5_2);
  nand NAND2_3889(II19717,WX5812,II19716);
  nand NAND2_3890(II19718,CRC_OUT_5_2,II19716);
  nand NAND2_3891(WX6432,II19717,II19718);
  nand NAND2_3892(II19723,WX5813,CRC_OUT_5_1);
  nand NAND2_3893(II19724,WX5813,II19723);
  nand NAND2_3894(II19725,CRC_OUT_5_1,II19723);
  nand NAND2_3895(WX6433,II19724,II19725);
  nand NAND2_3896(II19730,WX5814,CRC_OUT_5_0);
  nand NAND2_3897(II19731,WX5814,II19730);
  nand NAND2_3898(II19732,CRC_OUT_5_0,II19730);
  nand NAND2_3899(WX6434,II19731,II19732);
  nand NAND2_3900(II22013,WX7466,WX7110);
  nand NAND2_3901(II22014,WX7466,II22013);
  nand NAND2_3902(II22015,WX7110,II22013);
  nand NAND2_3903(II22012,II22014,II22015);
  nand NAND2_3904(II22020,WX7174,II22012);
  nand NAND2_3905(II22021,WX7174,II22020);
  nand NAND2_3906(II22022,II22012,II22020);
  nand NAND2_3907(II22011,II22021,II22022);
  nand NAND2_3908(II22028,WX7238,WX7302);
  nand NAND2_3909(II22029,WX7238,II22028);
  nand NAND2_3910(II22030,WX7302,II22028);
  nand NAND2_3911(II22027,II22029,II22030);
  nand NAND2_3912(II22035,II22011,II22027);
  nand NAND2_3913(II22036,II22011,II22035);
  nand NAND2_3914(II22037,II22027,II22035);
  nand NAND2_3915(WX7365,II22036,II22037);
  nand NAND2_3916(II22044,WX7466,WX7112);
  nand NAND2_3917(II22045,WX7466,II22044);
  nand NAND2_3918(II22046,WX7112,II22044);
  nand NAND2_3919(II22043,II22045,II22046);
  nand NAND2_3920(II22051,WX7176,II22043);
  nand NAND2_3921(II22052,WX7176,II22051);
  nand NAND2_3922(II22053,II22043,II22051);
  nand NAND2_3923(II22042,II22052,II22053);
  nand NAND2_3924(II22059,WX7240,WX7304);
  nand NAND2_3925(II22060,WX7240,II22059);
  nand NAND2_3926(II22061,WX7304,II22059);
  nand NAND2_3927(II22058,II22060,II22061);
  nand NAND2_3928(II22066,II22042,II22058);
  nand NAND2_3929(II22067,II22042,II22066);
  nand NAND2_3930(II22068,II22058,II22066);
  nand NAND2_3931(WX7366,II22067,II22068);
  nand NAND2_3932(II22075,WX7466,WX7114);
  nand NAND2_3933(II22076,WX7466,II22075);
  nand NAND2_3934(II22077,WX7114,II22075);
  nand NAND2_3935(II22074,II22076,II22077);
  nand NAND2_3936(II22082,WX7178,II22074);
  nand NAND2_3937(II22083,WX7178,II22082);
  nand NAND2_3938(II22084,II22074,II22082);
  nand NAND2_3939(II22073,II22083,II22084);
  nand NAND2_3940(II22090,WX7242,WX7306);
  nand NAND2_3941(II22091,WX7242,II22090);
  nand NAND2_3942(II22092,WX7306,II22090);
  nand NAND2_3943(II22089,II22091,II22092);
  nand NAND2_3944(II22097,II22073,II22089);
  nand NAND2_3945(II22098,II22073,II22097);
  nand NAND2_3946(II22099,II22089,II22097);
  nand NAND2_3947(WX7367,II22098,II22099);
  nand NAND2_3948(II22106,WX7466,WX7116);
  nand NAND2_3949(II22107,WX7466,II22106);
  nand NAND2_3950(II22108,WX7116,II22106);
  nand NAND2_3951(II22105,II22107,II22108);
  nand NAND2_3952(II22113,WX7180,II22105);
  nand NAND2_3953(II22114,WX7180,II22113);
  nand NAND2_3954(II22115,II22105,II22113);
  nand NAND2_3955(II22104,II22114,II22115);
  nand NAND2_3956(II22121,WX7244,WX7308);
  nand NAND2_3957(II22122,WX7244,II22121);
  nand NAND2_3958(II22123,WX7308,II22121);
  nand NAND2_3959(II22120,II22122,II22123);
  nand NAND2_3960(II22128,II22104,II22120);
  nand NAND2_3961(II22129,II22104,II22128);
  nand NAND2_3962(II22130,II22120,II22128);
  nand NAND2_3963(WX7368,II22129,II22130);
  nand NAND2_3964(II22137,WX7466,WX7118);
  nand NAND2_3965(II22138,WX7466,II22137);
  nand NAND2_3966(II22139,WX7118,II22137);
  nand NAND2_3967(II22136,II22138,II22139);
  nand NAND2_3968(II22144,WX7182,II22136);
  nand NAND2_3969(II22145,WX7182,II22144);
  nand NAND2_3970(II22146,II22136,II22144);
  nand NAND2_3971(II22135,II22145,II22146);
  nand NAND2_3972(II22152,WX7246,WX7310);
  nand NAND2_3973(II22153,WX7246,II22152);
  nand NAND2_3974(II22154,WX7310,II22152);
  nand NAND2_3975(II22151,II22153,II22154);
  nand NAND2_3976(II22159,II22135,II22151);
  nand NAND2_3977(II22160,II22135,II22159);
  nand NAND2_3978(II22161,II22151,II22159);
  nand NAND2_3979(WX7369,II22160,II22161);
  nand NAND2_3980(II22168,WX7466,WX7120);
  nand NAND2_3981(II22169,WX7466,II22168);
  nand NAND2_3982(II22170,WX7120,II22168);
  nand NAND2_3983(II22167,II22169,II22170);
  nand NAND2_3984(II22175,WX7184,II22167);
  nand NAND2_3985(II22176,WX7184,II22175);
  nand NAND2_3986(II22177,II22167,II22175);
  nand NAND2_3987(II22166,II22176,II22177);
  nand NAND2_3988(II22183,WX7248,WX7312);
  nand NAND2_3989(II22184,WX7248,II22183);
  nand NAND2_3990(II22185,WX7312,II22183);
  nand NAND2_3991(II22182,II22184,II22185);
  nand NAND2_3992(II22190,II22166,II22182);
  nand NAND2_3993(II22191,II22166,II22190);
  nand NAND2_3994(II22192,II22182,II22190);
  nand NAND2_3995(WX7370,II22191,II22192);
  nand NAND2_3996(II22199,WX7466,WX7122);
  nand NAND2_3997(II22200,WX7466,II22199);
  nand NAND2_3998(II22201,WX7122,II22199);
  nand NAND2_3999(II22198,II22200,II22201);
  nand NAND2_4000(II22206,WX7186,II22198);
  nand NAND2_4001(II22207,WX7186,II22206);
  nand NAND2_4002(II22208,II22198,II22206);
  nand NAND2_4003(II22197,II22207,II22208);
  nand NAND2_4004(II22214,WX7250,WX7314);
  nand NAND2_4005(II22215,WX7250,II22214);
  nand NAND2_4006(II22216,WX7314,II22214);
  nand NAND2_4007(II22213,II22215,II22216);
  nand NAND2_4008(II22221,II22197,II22213);
  nand NAND2_4009(II22222,II22197,II22221);
  nand NAND2_4010(II22223,II22213,II22221);
  nand NAND2_4011(WX7371,II22222,II22223);
  nand NAND2_4012(II22230,WX7466,WX7124);
  nand NAND2_4013(II22231,WX7466,II22230);
  nand NAND2_4014(II22232,WX7124,II22230);
  nand NAND2_4015(II22229,II22231,II22232);
  nand NAND2_4016(II22237,WX7188,II22229);
  nand NAND2_4017(II22238,WX7188,II22237);
  nand NAND2_4018(II22239,II22229,II22237);
  nand NAND2_4019(II22228,II22238,II22239);
  nand NAND2_4020(II22245,WX7252,WX7316);
  nand NAND2_4021(II22246,WX7252,II22245);
  nand NAND2_4022(II22247,WX7316,II22245);
  nand NAND2_4023(II22244,II22246,II22247);
  nand NAND2_4024(II22252,II22228,II22244);
  nand NAND2_4025(II22253,II22228,II22252);
  nand NAND2_4026(II22254,II22244,II22252);
  nand NAND2_4027(WX7372,II22253,II22254);
  nand NAND2_4028(II22261,WX7466,WX7126);
  nand NAND2_4029(II22262,WX7466,II22261);
  nand NAND2_4030(II22263,WX7126,II22261);
  nand NAND2_4031(II22260,II22262,II22263);
  nand NAND2_4032(II22268,WX7190,II22260);
  nand NAND2_4033(II22269,WX7190,II22268);
  nand NAND2_4034(II22270,II22260,II22268);
  nand NAND2_4035(II22259,II22269,II22270);
  nand NAND2_4036(II22276,WX7254,WX7318);
  nand NAND2_4037(II22277,WX7254,II22276);
  nand NAND2_4038(II22278,WX7318,II22276);
  nand NAND2_4039(II22275,II22277,II22278);
  nand NAND2_4040(II22283,II22259,II22275);
  nand NAND2_4041(II22284,II22259,II22283);
  nand NAND2_4042(II22285,II22275,II22283);
  nand NAND2_4043(WX7373,II22284,II22285);
  nand NAND2_4044(II22292,WX7466,WX7128);
  nand NAND2_4045(II22293,WX7466,II22292);
  nand NAND2_4046(II22294,WX7128,II22292);
  nand NAND2_4047(II22291,II22293,II22294);
  nand NAND2_4048(II22299,WX7192,II22291);
  nand NAND2_4049(II22300,WX7192,II22299);
  nand NAND2_4050(II22301,II22291,II22299);
  nand NAND2_4051(II22290,II22300,II22301);
  nand NAND2_4052(II22307,WX7256,WX7320);
  nand NAND2_4053(II22308,WX7256,II22307);
  nand NAND2_4054(II22309,WX7320,II22307);
  nand NAND2_4055(II22306,II22308,II22309);
  nand NAND2_4056(II22314,II22290,II22306);
  nand NAND2_4057(II22315,II22290,II22314);
  nand NAND2_4058(II22316,II22306,II22314);
  nand NAND2_4059(WX7374,II22315,II22316);
  nand NAND2_4060(II22323,WX7466,WX7130);
  nand NAND2_4061(II22324,WX7466,II22323);
  nand NAND2_4062(II22325,WX7130,II22323);
  nand NAND2_4063(II22322,II22324,II22325);
  nand NAND2_4064(II22330,WX7194,II22322);
  nand NAND2_4065(II22331,WX7194,II22330);
  nand NAND2_4066(II22332,II22322,II22330);
  nand NAND2_4067(II22321,II22331,II22332);
  nand NAND2_4068(II22338,WX7258,WX7322);
  nand NAND2_4069(II22339,WX7258,II22338);
  nand NAND2_4070(II22340,WX7322,II22338);
  nand NAND2_4071(II22337,II22339,II22340);
  nand NAND2_4072(II22345,II22321,II22337);
  nand NAND2_4073(II22346,II22321,II22345);
  nand NAND2_4074(II22347,II22337,II22345);
  nand NAND2_4075(WX7375,II22346,II22347);
  nand NAND2_4076(II22354,WX7466,WX7132);
  nand NAND2_4077(II22355,WX7466,II22354);
  nand NAND2_4078(II22356,WX7132,II22354);
  nand NAND2_4079(II22353,II22355,II22356);
  nand NAND2_4080(II22361,WX7196,II22353);
  nand NAND2_4081(II22362,WX7196,II22361);
  nand NAND2_4082(II22363,II22353,II22361);
  nand NAND2_4083(II22352,II22362,II22363);
  nand NAND2_4084(II22369,WX7260,WX7324);
  nand NAND2_4085(II22370,WX7260,II22369);
  nand NAND2_4086(II22371,WX7324,II22369);
  nand NAND2_4087(II22368,II22370,II22371);
  nand NAND2_4088(II22376,II22352,II22368);
  nand NAND2_4089(II22377,II22352,II22376);
  nand NAND2_4090(II22378,II22368,II22376);
  nand NAND2_4091(WX7376,II22377,II22378);
  nand NAND2_4092(II22385,WX7466,WX7134);
  nand NAND2_4093(II22386,WX7466,II22385);
  nand NAND2_4094(II22387,WX7134,II22385);
  nand NAND2_4095(II22384,II22386,II22387);
  nand NAND2_4096(II22392,WX7198,II22384);
  nand NAND2_4097(II22393,WX7198,II22392);
  nand NAND2_4098(II22394,II22384,II22392);
  nand NAND2_4099(II22383,II22393,II22394);
  nand NAND2_4100(II22400,WX7262,WX7326);
  nand NAND2_4101(II22401,WX7262,II22400);
  nand NAND2_4102(II22402,WX7326,II22400);
  nand NAND2_4103(II22399,II22401,II22402);
  nand NAND2_4104(II22407,II22383,II22399);
  nand NAND2_4105(II22408,II22383,II22407);
  nand NAND2_4106(II22409,II22399,II22407);
  nand NAND2_4107(WX7377,II22408,II22409);
  nand NAND2_4108(II22416,WX7466,WX7136);
  nand NAND2_4109(II22417,WX7466,II22416);
  nand NAND2_4110(II22418,WX7136,II22416);
  nand NAND2_4111(II22415,II22417,II22418);
  nand NAND2_4112(II22423,WX7200,II22415);
  nand NAND2_4113(II22424,WX7200,II22423);
  nand NAND2_4114(II22425,II22415,II22423);
  nand NAND2_4115(II22414,II22424,II22425);
  nand NAND2_4116(II22431,WX7264,WX7328);
  nand NAND2_4117(II22432,WX7264,II22431);
  nand NAND2_4118(II22433,WX7328,II22431);
  nand NAND2_4119(II22430,II22432,II22433);
  nand NAND2_4120(II22438,II22414,II22430);
  nand NAND2_4121(II22439,II22414,II22438);
  nand NAND2_4122(II22440,II22430,II22438);
  nand NAND2_4123(WX7378,II22439,II22440);
  nand NAND2_4124(II22447,WX7466,WX7138);
  nand NAND2_4125(II22448,WX7466,II22447);
  nand NAND2_4126(II22449,WX7138,II22447);
  nand NAND2_4127(II22446,II22448,II22449);
  nand NAND2_4128(II22454,WX7202,II22446);
  nand NAND2_4129(II22455,WX7202,II22454);
  nand NAND2_4130(II22456,II22446,II22454);
  nand NAND2_4131(II22445,II22455,II22456);
  nand NAND2_4132(II22462,WX7266,WX7330);
  nand NAND2_4133(II22463,WX7266,II22462);
  nand NAND2_4134(II22464,WX7330,II22462);
  nand NAND2_4135(II22461,II22463,II22464);
  nand NAND2_4136(II22469,II22445,II22461);
  nand NAND2_4137(II22470,II22445,II22469);
  nand NAND2_4138(II22471,II22461,II22469);
  nand NAND2_4139(WX7379,II22470,II22471);
  nand NAND2_4140(II22478,WX7466,WX7140);
  nand NAND2_4141(II22479,WX7466,II22478);
  nand NAND2_4142(II22480,WX7140,II22478);
  nand NAND2_4143(II22477,II22479,II22480);
  nand NAND2_4144(II22485,WX7204,II22477);
  nand NAND2_4145(II22486,WX7204,II22485);
  nand NAND2_4146(II22487,II22477,II22485);
  nand NAND2_4147(II22476,II22486,II22487);
  nand NAND2_4148(II22493,WX7268,WX7332);
  nand NAND2_4149(II22494,WX7268,II22493);
  nand NAND2_4150(II22495,WX7332,II22493);
  nand NAND2_4151(II22492,II22494,II22495);
  nand NAND2_4152(II22500,II22476,II22492);
  nand NAND2_4153(II22501,II22476,II22500);
  nand NAND2_4154(II22502,II22492,II22500);
  nand NAND2_4155(WX7380,II22501,II22502);
  nand NAND2_4156(II22509,WX7467,WX7142);
  nand NAND2_4157(II22510,WX7467,II22509);
  nand NAND2_4158(II22511,WX7142,II22509);
  nand NAND2_4159(II22508,II22510,II22511);
  nand NAND2_4160(II22516,WX7206,II22508);
  nand NAND2_4161(II22517,WX7206,II22516);
  nand NAND2_4162(II22518,II22508,II22516);
  nand NAND2_4163(II22507,II22517,II22518);
  nand NAND2_4164(II22524,WX7270,WX7334);
  nand NAND2_4165(II22525,WX7270,II22524);
  nand NAND2_4166(II22526,WX7334,II22524);
  nand NAND2_4167(II22523,II22525,II22526);
  nand NAND2_4168(II22531,II22507,II22523);
  nand NAND2_4169(II22532,II22507,II22531);
  nand NAND2_4170(II22533,II22523,II22531);
  nand NAND2_4171(WX7381,II22532,II22533);
  nand NAND2_4172(II22540,WX7467,WX7144);
  nand NAND2_4173(II22541,WX7467,II22540);
  nand NAND2_4174(II22542,WX7144,II22540);
  nand NAND2_4175(II22539,II22541,II22542);
  nand NAND2_4176(II22547,WX7208,II22539);
  nand NAND2_4177(II22548,WX7208,II22547);
  nand NAND2_4178(II22549,II22539,II22547);
  nand NAND2_4179(II22538,II22548,II22549);
  nand NAND2_4180(II22555,WX7272,WX7336);
  nand NAND2_4181(II22556,WX7272,II22555);
  nand NAND2_4182(II22557,WX7336,II22555);
  nand NAND2_4183(II22554,II22556,II22557);
  nand NAND2_4184(II22562,II22538,II22554);
  nand NAND2_4185(II22563,II22538,II22562);
  nand NAND2_4186(II22564,II22554,II22562);
  nand NAND2_4187(WX7382,II22563,II22564);
  nand NAND2_4188(II22571,WX7467,WX7146);
  nand NAND2_4189(II22572,WX7467,II22571);
  nand NAND2_4190(II22573,WX7146,II22571);
  nand NAND2_4191(II22570,II22572,II22573);
  nand NAND2_4192(II22578,WX7210,II22570);
  nand NAND2_4193(II22579,WX7210,II22578);
  nand NAND2_4194(II22580,II22570,II22578);
  nand NAND2_4195(II22569,II22579,II22580);
  nand NAND2_4196(II22586,WX7274,WX7338);
  nand NAND2_4197(II22587,WX7274,II22586);
  nand NAND2_4198(II22588,WX7338,II22586);
  nand NAND2_4199(II22585,II22587,II22588);
  nand NAND2_4200(II22593,II22569,II22585);
  nand NAND2_4201(II22594,II22569,II22593);
  nand NAND2_4202(II22595,II22585,II22593);
  nand NAND2_4203(WX7383,II22594,II22595);
  nand NAND2_4204(II22602,WX7467,WX7148);
  nand NAND2_4205(II22603,WX7467,II22602);
  nand NAND2_4206(II22604,WX7148,II22602);
  nand NAND2_4207(II22601,II22603,II22604);
  nand NAND2_4208(II22609,WX7212,II22601);
  nand NAND2_4209(II22610,WX7212,II22609);
  nand NAND2_4210(II22611,II22601,II22609);
  nand NAND2_4211(II22600,II22610,II22611);
  nand NAND2_4212(II22617,WX7276,WX7340);
  nand NAND2_4213(II22618,WX7276,II22617);
  nand NAND2_4214(II22619,WX7340,II22617);
  nand NAND2_4215(II22616,II22618,II22619);
  nand NAND2_4216(II22624,II22600,II22616);
  nand NAND2_4217(II22625,II22600,II22624);
  nand NAND2_4218(II22626,II22616,II22624);
  nand NAND2_4219(WX7384,II22625,II22626);
  nand NAND2_4220(II22633,WX7467,WX7150);
  nand NAND2_4221(II22634,WX7467,II22633);
  nand NAND2_4222(II22635,WX7150,II22633);
  nand NAND2_4223(II22632,II22634,II22635);
  nand NAND2_4224(II22640,WX7214,II22632);
  nand NAND2_4225(II22641,WX7214,II22640);
  nand NAND2_4226(II22642,II22632,II22640);
  nand NAND2_4227(II22631,II22641,II22642);
  nand NAND2_4228(II22648,WX7278,WX7342);
  nand NAND2_4229(II22649,WX7278,II22648);
  nand NAND2_4230(II22650,WX7342,II22648);
  nand NAND2_4231(II22647,II22649,II22650);
  nand NAND2_4232(II22655,II22631,II22647);
  nand NAND2_4233(II22656,II22631,II22655);
  nand NAND2_4234(II22657,II22647,II22655);
  nand NAND2_4235(WX7385,II22656,II22657);
  nand NAND2_4236(II22664,WX7467,WX7152);
  nand NAND2_4237(II22665,WX7467,II22664);
  nand NAND2_4238(II22666,WX7152,II22664);
  nand NAND2_4239(II22663,II22665,II22666);
  nand NAND2_4240(II22671,WX7216,II22663);
  nand NAND2_4241(II22672,WX7216,II22671);
  nand NAND2_4242(II22673,II22663,II22671);
  nand NAND2_4243(II22662,II22672,II22673);
  nand NAND2_4244(II22679,WX7280,WX7344);
  nand NAND2_4245(II22680,WX7280,II22679);
  nand NAND2_4246(II22681,WX7344,II22679);
  nand NAND2_4247(II22678,II22680,II22681);
  nand NAND2_4248(II22686,II22662,II22678);
  nand NAND2_4249(II22687,II22662,II22686);
  nand NAND2_4250(II22688,II22678,II22686);
  nand NAND2_4251(WX7386,II22687,II22688);
  nand NAND2_4252(II22695,WX7467,WX7154);
  nand NAND2_4253(II22696,WX7467,II22695);
  nand NAND2_4254(II22697,WX7154,II22695);
  nand NAND2_4255(II22694,II22696,II22697);
  nand NAND2_4256(II22702,WX7218,II22694);
  nand NAND2_4257(II22703,WX7218,II22702);
  nand NAND2_4258(II22704,II22694,II22702);
  nand NAND2_4259(II22693,II22703,II22704);
  nand NAND2_4260(II22710,WX7282,WX7346);
  nand NAND2_4261(II22711,WX7282,II22710);
  nand NAND2_4262(II22712,WX7346,II22710);
  nand NAND2_4263(II22709,II22711,II22712);
  nand NAND2_4264(II22717,II22693,II22709);
  nand NAND2_4265(II22718,II22693,II22717);
  nand NAND2_4266(II22719,II22709,II22717);
  nand NAND2_4267(WX7387,II22718,II22719);
  nand NAND2_4268(II22726,WX7467,WX7156);
  nand NAND2_4269(II22727,WX7467,II22726);
  nand NAND2_4270(II22728,WX7156,II22726);
  nand NAND2_4271(II22725,II22727,II22728);
  nand NAND2_4272(II22733,WX7220,II22725);
  nand NAND2_4273(II22734,WX7220,II22733);
  nand NAND2_4274(II22735,II22725,II22733);
  nand NAND2_4275(II22724,II22734,II22735);
  nand NAND2_4276(II22741,WX7284,WX7348);
  nand NAND2_4277(II22742,WX7284,II22741);
  nand NAND2_4278(II22743,WX7348,II22741);
  nand NAND2_4279(II22740,II22742,II22743);
  nand NAND2_4280(II22748,II22724,II22740);
  nand NAND2_4281(II22749,II22724,II22748);
  nand NAND2_4282(II22750,II22740,II22748);
  nand NAND2_4283(WX7388,II22749,II22750);
  nand NAND2_4284(II22757,WX7467,WX7158);
  nand NAND2_4285(II22758,WX7467,II22757);
  nand NAND2_4286(II22759,WX7158,II22757);
  nand NAND2_4287(II22756,II22758,II22759);
  nand NAND2_4288(II22764,WX7222,II22756);
  nand NAND2_4289(II22765,WX7222,II22764);
  nand NAND2_4290(II22766,II22756,II22764);
  nand NAND2_4291(II22755,II22765,II22766);
  nand NAND2_4292(II22772,WX7286,WX7350);
  nand NAND2_4293(II22773,WX7286,II22772);
  nand NAND2_4294(II22774,WX7350,II22772);
  nand NAND2_4295(II22771,II22773,II22774);
  nand NAND2_4296(II22779,II22755,II22771);
  nand NAND2_4297(II22780,II22755,II22779);
  nand NAND2_4298(II22781,II22771,II22779);
  nand NAND2_4299(WX7389,II22780,II22781);
  nand NAND2_4300(II22788,WX7467,WX7160);
  nand NAND2_4301(II22789,WX7467,II22788);
  nand NAND2_4302(II22790,WX7160,II22788);
  nand NAND2_4303(II22787,II22789,II22790);
  nand NAND2_4304(II22795,WX7224,II22787);
  nand NAND2_4305(II22796,WX7224,II22795);
  nand NAND2_4306(II22797,II22787,II22795);
  nand NAND2_4307(II22786,II22796,II22797);
  nand NAND2_4308(II22803,WX7288,WX7352);
  nand NAND2_4309(II22804,WX7288,II22803);
  nand NAND2_4310(II22805,WX7352,II22803);
  nand NAND2_4311(II22802,II22804,II22805);
  nand NAND2_4312(II22810,II22786,II22802);
  nand NAND2_4313(II22811,II22786,II22810);
  nand NAND2_4314(II22812,II22802,II22810);
  nand NAND2_4315(WX7390,II22811,II22812);
  nand NAND2_4316(II22819,WX7467,WX7162);
  nand NAND2_4317(II22820,WX7467,II22819);
  nand NAND2_4318(II22821,WX7162,II22819);
  nand NAND2_4319(II22818,II22820,II22821);
  nand NAND2_4320(II22826,WX7226,II22818);
  nand NAND2_4321(II22827,WX7226,II22826);
  nand NAND2_4322(II22828,II22818,II22826);
  nand NAND2_4323(II22817,II22827,II22828);
  nand NAND2_4324(II22834,WX7290,WX7354);
  nand NAND2_4325(II22835,WX7290,II22834);
  nand NAND2_4326(II22836,WX7354,II22834);
  nand NAND2_4327(II22833,II22835,II22836);
  nand NAND2_4328(II22841,II22817,II22833);
  nand NAND2_4329(II22842,II22817,II22841);
  nand NAND2_4330(II22843,II22833,II22841);
  nand NAND2_4331(WX7391,II22842,II22843);
  nand NAND2_4332(II22850,WX7467,WX7164);
  nand NAND2_4333(II22851,WX7467,II22850);
  nand NAND2_4334(II22852,WX7164,II22850);
  nand NAND2_4335(II22849,II22851,II22852);
  nand NAND2_4336(II22857,WX7228,II22849);
  nand NAND2_4337(II22858,WX7228,II22857);
  nand NAND2_4338(II22859,II22849,II22857);
  nand NAND2_4339(II22848,II22858,II22859);
  nand NAND2_4340(II22865,WX7292,WX7356);
  nand NAND2_4341(II22866,WX7292,II22865);
  nand NAND2_4342(II22867,WX7356,II22865);
  nand NAND2_4343(II22864,II22866,II22867);
  nand NAND2_4344(II22872,II22848,II22864);
  nand NAND2_4345(II22873,II22848,II22872);
  nand NAND2_4346(II22874,II22864,II22872);
  nand NAND2_4347(WX7392,II22873,II22874);
  nand NAND2_4348(II22881,WX7467,WX7166);
  nand NAND2_4349(II22882,WX7467,II22881);
  nand NAND2_4350(II22883,WX7166,II22881);
  nand NAND2_4351(II22880,II22882,II22883);
  nand NAND2_4352(II22888,WX7230,II22880);
  nand NAND2_4353(II22889,WX7230,II22888);
  nand NAND2_4354(II22890,II22880,II22888);
  nand NAND2_4355(II22879,II22889,II22890);
  nand NAND2_4356(II22896,WX7294,WX7358);
  nand NAND2_4357(II22897,WX7294,II22896);
  nand NAND2_4358(II22898,WX7358,II22896);
  nand NAND2_4359(II22895,II22897,II22898);
  nand NAND2_4360(II22903,II22879,II22895);
  nand NAND2_4361(II22904,II22879,II22903);
  nand NAND2_4362(II22905,II22895,II22903);
  nand NAND2_4363(WX7393,II22904,II22905);
  nand NAND2_4364(II22912,WX7467,WX7168);
  nand NAND2_4365(II22913,WX7467,II22912);
  nand NAND2_4366(II22914,WX7168,II22912);
  nand NAND2_4367(II22911,II22913,II22914);
  nand NAND2_4368(II22919,WX7232,II22911);
  nand NAND2_4369(II22920,WX7232,II22919);
  nand NAND2_4370(II22921,II22911,II22919);
  nand NAND2_4371(II22910,II22920,II22921);
  nand NAND2_4372(II22927,WX7296,WX7360);
  nand NAND2_4373(II22928,WX7296,II22927);
  nand NAND2_4374(II22929,WX7360,II22927);
  nand NAND2_4375(II22926,II22928,II22929);
  nand NAND2_4376(II22934,II22910,II22926);
  nand NAND2_4377(II22935,II22910,II22934);
  nand NAND2_4378(II22936,II22926,II22934);
  nand NAND2_4379(WX7394,II22935,II22936);
  nand NAND2_4380(II22943,WX7467,WX7170);
  nand NAND2_4381(II22944,WX7467,II22943);
  nand NAND2_4382(II22945,WX7170,II22943);
  nand NAND2_4383(II22942,II22944,II22945);
  nand NAND2_4384(II22950,WX7234,II22942);
  nand NAND2_4385(II22951,WX7234,II22950);
  nand NAND2_4386(II22952,II22942,II22950);
  nand NAND2_4387(II22941,II22951,II22952);
  nand NAND2_4388(II22958,WX7298,WX7362);
  nand NAND2_4389(II22959,WX7298,II22958);
  nand NAND2_4390(II22960,WX7362,II22958);
  nand NAND2_4391(II22957,II22959,II22960);
  nand NAND2_4392(II22965,II22941,II22957);
  nand NAND2_4393(II22966,II22941,II22965);
  nand NAND2_4394(II22967,II22957,II22965);
  nand NAND2_4395(WX7395,II22966,II22967);
  nand NAND2_4396(II22974,WX7467,WX7172);
  nand NAND2_4397(II22975,WX7467,II22974);
  nand NAND2_4398(II22976,WX7172,II22974);
  nand NAND2_4399(II22973,II22975,II22976);
  nand NAND2_4400(II22981,WX7236,II22973);
  nand NAND2_4401(II22982,WX7236,II22981);
  nand NAND2_4402(II22983,II22973,II22981);
  nand NAND2_4403(II22972,II22982,II22983);
  nand NAND2_4404(II22989,WX7300,WX7364);
  nand NAND2_4405(II22990,WX7300,II22989);
  nand NAND2_4406(II22991,WX7364,II22989);
  nand NAND2_4407(II22988,II22990,II22991);
  nand NAND2_4408(II22996,II22972,II22988);
  nand NAND2_4409(II22997,II22972,II22996);
  nand NAND2_4410(II22998,II22988,II22996);
  nand NAND2_4411(WX7396,II22997,II22998);
  nand NAND2_4412(II23077,WX7045,WX6950);
  nand NAND2_4413(II23078,WX7045,II23077);
  nand NAND2_4414(II23079,WX6950,II23077);
  nand NAND2_4415(WX7471,II23078,II23079);
  nand NAND2_4416(II23090,WX7046,WX6952);
  nand NAND2_4417(II23091,WX7046,II23090);
  nand NAND2_4418(II23092,WX6952,II23090);
  nand NAND2_4419(WX7478,II23091,II23092);
  nand NAND2_4420(II23103,WX7047,WX6954);
  nand NAND2_4421(II23104,WX7047,II23103);
  nand NAND2_4422(II23105,WX6954,II23103);
  nand NAND2_4423(WX7485,II23104,II23105);
  nand NAND2_4424(II23116,WX7048,WX6956);
  nand NAND2_4425(II23117,WX7048,II23116);
  nand NAND2_4426(II23118,WX6956,II23116);
  nand NAND2_4427(WX7492,II23117,II23118);
  nand NAND2_4428(II23129,WX7049,WX6958);
  nand NAND2_4429(II23130,WX7049,II23129);
  nand NAND2_4430(II23131,WX6958,II23129);
  nand NAND2_4431(WX7499,II23130,II23131);
  nand NAND2_4432(II23142,WX7050,WX6960);
  nand NAND2_4433(II23143,WX7050,II23142);
  nand NAND2_4434(II23144,WX6960,II23142);
  nand NAND2_4435(WX7506,II23143,II23144);
  nand NAND2_4436(II23155,WX7051,WX6962);
  nand NAND2_4437(II23156,WX7051,II23155);
  nand NAND2_4438(II23157,WX6962,II23155);
  nand NAND2_4439(WX7513,II23156,II23157);
  nand NAND2_4440(II23168,WX7052,WX6964);
  nand NAND2_4441(II23169,WX7052,II23168);
  nand NAND2_4442(II23170,WX6964,II23168);
  nand NAND2_4443(WX7520,II23169,II23170);
  nand NAND2_4444(II23181,WX7053,WX6966);
  nand NAND2_4445(II23182,WX7053,II23181);
  nand NAND2_4446(II23183,WX6966,II23181);
  nand NAND2_4447(WX7527,II23182,II23183);
  nand NAND2_4448(II23194,WX7054,WX6968);
  nand NAND2_4449(II23195,WX7054,II23194);
  nand NAND2_4450(II23196,WX6968,II23194);
  nand NAND2_4451(WX7534,II23195,II23196);
  nand NAND2_4452(II23207,WX7055,WX6970);
  nand NAND2_4453(II23208,WX7055,II23207);
  nand NAND2_4454(II23209,WX6970,II23207);
  nand NAND2_4455(WX7541,II23208,II23209);
  nand NAND2_4456(II23220,WX7056,WX6972);
  nand NAND2_4457(II23221,WX7056,II23220);
  nand NAND2_4458(II23222,WX6972,II23220);
  nand NAND2_4459(WX7548,II23221,II23222);
  nand NAND2_4460(II23233,WX7057,WX6974);
  nand NAND2_4461(II23234,WX7057,II23233);
  nand NAND2_4462(II23235,WX6974,II23233);
  nand NAND2_4463(WX7555,II23234,II23235);
  nand NAND2_4464(II23246,WX7058,WX6976);
  nand NAND2_4465(II23247,WX7058,II23246);
  nand NAND2_4466(II23248,WX6976,II23246);
  nand NAND2_4467(WX7562,II23247,II23248);
  nand NAND2_4468(II23259,WX7059,WX6978);
  nand NAND2_4469(II23260,WX7059,II23259);
  nand NAND2_4470(II23261,WX6978,II23259);
  nand NAND2_4471(WX7569,II23260,II23261);
  nand NAND2_4472(II23272,WX7060,WX6980);
  nand NAND2_4473(II23273,WX7060,II23272);
  nand NAND2_4474(II23274,WX6980,II23272);
  nand NAND2_4475(WX7576,II23273,II23274);
  nand NAND2_4476(II23285,WX7061,WX6982);
  nand NAND2_4477(II23286,WX7061,II23285);
  nand NAND2_4478(II23287,WX6982,II23285);
  nand NAND2_4479(WX7583,II23286,II23287);
  nand NAND2_4480(II23298,WX7062,WX6984);
  nand NAND2_4481(II23299,WX7062,II23298);
  nand NAND2_4482(II23300,WX6984,II23298);
  nand NAND2_4483(WX7590,II23299,II23300);
  nand NAND2_4484(II23311,WX7063,WX6986);
  nand NAND2_4485(II23312,WX7063,II23311);
  nand NAND2_4486(II23313,WX6986,II23311);
  nand NAND2_4487(WX7597,II23312,II23313);
  nand NAND2_4488(II23324,WX7064,WX6988);
  nand NAND2_4489(II23325,WX7064,II23324);
  nand NAND2_4490(II23326,WX6988,II23324);
  nand NAND2_4491(WX7604,II23325,II23326);
  nand NAND2_4492(II23337,WX7065,WX6990);
  nand NAND2_4493(II23338,WX7065,II23337);
  nand NAND2_4494(II23339,WX6990,II23337);
  nand NAND2_4495(WX7611,II23338,II23339);
  nand NAND2_4496(II23350,WX7066,WX6992);
  nand NAND2_4497(II23351,WX7066,II23350);
  nand NAND2_4498(II23352,WX6992,II23350);
  nand NAND2_4499(WX7618,II23351,II23352);
  nand NAND2_4500(II23363,WX7067,WX6994);
  nand NAND2_4501(II23364,WX7067,II23363);
  nand NAND2_4502(II23365,WX6994,II23363);
  nand NAND2_4503(WX7625,II23364,II23365);
  nand NAND2_4504(II23376,WX7068,WX6996);
  nand NAND2_4505(II23377,WX7068,II23376);
  nand NAND2_4506(II23378,WX6996,II23376);
  nand NAND2_4507(WX7632,II23377,II23378);
  nand NAND2_4508(II23389,WX7069,WX6998);
  nand NAND2_4509(II23390,WX7069,II23389);
  nand NAND2_4510(II23391,WX6998,II23389);
  nand NAND2_4511(WX7639,II23390,II23391);
  nand NAND2_4512(II23402,WX7070,WX7000);
  nand NAND2_4513(II23403,WX7070,II23402);
  nand NAND2_4514(II23404,WX7000,II23402);
  nand NAND2_4515(WX7646,II23403,II23404);
  nand NAND2_4516(II23415,WX7071,WX7002);
  nand NAND2_4517(II23416,WX7071,II23415);
  nand NAND2_4518(II23417,WX7002,II23415);
  nand NAND2_4519(WX7653,II23416,II23417);
  nand NAND2_4520(II23428,WX7072,WX7004);
  nand NAND2_4521(II23429,WX7072,II23428);
  nand NAND2_4522(II23430,WX7004,II23428);
  nand NAND2_4523(WX7660,II23429,II23430);
  nand NAND2_4524(II23441,WX7073,WX7006);
  nand NAND2_4525(II23442,WX7073,II23441);
  nand NAND2_4526(II23443,WX7006,II23441);
  nand NAND2_4527(WX7667,II23442,II23443);
  nand NAND2_4528(II23454,WX7074,WX7008);
  nand NAND2_4529(II23455,WX7074,II23454);
  nand NAND2_4530(II23456,WX7008,II23454);
  nand NAND2_4531(WX7674,II23455,II23456);
  nand NAND2_4532(II23467,WX7075,WX7010);
  nand NAND2_4533(II23468,WX7075,II23467);
  nand NAND2_4534(II23469,WX7010,II23467);
  nand NAND2_4535(WX7681,II23468,II23469);
  nand NAND2_4536(II23480,WX7076,WX7012);
  nand NAND2_4537(II23481,WX7076,II23480);
  nand NAND2_4538(II23482,WX7012,II23480);
  nand NAND2_4539(WX7688,II23481,II23482);
  nand NAND2_4540(II23495,WX7092,CRC_OUT_4_31);
  nand NAND2_4541(II23496,WX7092,II23495);
  nand NAND2_4542(II23497,CRC_OUT_4_31,II23495);
  nand NAND2_4543(II23494,II23496,II23497);
  nand NAND2_4544(II23502,CRC_OUT_4_15,II23494);
  nand NAND2_4545(II23503,CRC_OUT_4_15,II23502);
  nand NAND2_4546(II23504,II23494,II23502);
  nand NAND2_4547(WX7696,II23503,II23504);
  nand NAND2_4548(II23510,WX7097,CRC_OUT_4_31);
  nand NAND2_4549(II23511,WX7097,II23510);
  nand NAND2_4550(II23512,CRC_OUT_4_31,II23510);
  nand NAND2_4551(II23509,II23511,II23512);
  nand NAND2_4552(II23517,CRC_OUT_4_10,II23509);
  nand NAND2_4553(II23518,CRC_OUT_4_10,II23517);
  nand NAND2_4554(II23519,II23509,II23517);
  nand NAND2_4555(WX7697,II23518,II23519);
  nand NAND2_4556(II23525,WX7104,CRC_OUT_4_31);
  nand NAND2_4557(II23526,WX7104,II23525);
  nand NAND2_4558(II23527,CRC_OUT_4_31,II23525);
  nand NAND2_4559(II23524,II23526,II23527);
  nand NAND2_4560(II23532,CRC_OUT_4_3,II23524);
  nand NAND2_4561(II23533,CRC_OUT_4_3,II23532);
  nand NAND2_4562(II23534,II23524,II23532);
  nand NAND2_4563(WX7698,II23533,II23534);
  nand NAND2_4564(II23539,WX7108,CRC_OUT_4_31);
  nand NAND2_4565(II23540,WX7108,II23539);
  nand NAND2_4566(II23541,CRC_OUT_4_31,II23539);
  nand NAND2_4567(WX7699,II23540,II23541);
  nand NAND2_4568(II23546,WX7077,CRC_OUT_4_30);
  nand NAND2_4569(II23547,WX7077,II23546);
  nand NAND2_4570(II23548,CRC_OUT_4_30,II23546);
  nand NAND2_4571(WX7700,II23547,II23548);
  nand NAND2_4572(II23553,WX7078,CRC_OUT_4_29);
  nand NAND2_4573(II23554,WX7078,II23553);
  nand NAND2_4574(II23555,CRC_OUT_4_29,II23553);
  nand NAND2_4575(WX7701,II23554,II23555);
  nand NAND2_4576(II23560,WX7079,CRC_OUT_4_28);
  nand NAND2_4577(II23561,WX7079,II23560);
  nand NAND2_4578(II23562,CRC_OUT_4_28,II23560);
  nand NAND2_4579(WX7702,II23561,II23562);
  nand NAND2_4580(II23567,WX7080,CRC_OUT_4_27);
  nand NAND2_4581(II23568,WX7080,II23567);
  nand NAND2_4582(II23569,CRC_OUT_4_27,II23567);
  nand NAND2_4583(WX7703,II23568,II23569);
  nand NAND2_4584(II23574,WX7081,CRC_OUT_4_26);
  nand NAND2_4585(II23575,WX7081,II23574);
  nand NAND2_4586(II23576,CRC_OUT_4_26,II23574);
  nand NAND2_4587(WX7704,II23575,II23576);
  nand NAND2_4588(II23581,WX7082,CRC_OUT_4_25);
  nand NAND2_4589(II23582,WX7082,II23581);
  nand NAND2_4590(II23583,CRC_OUT_4_25,II23581);
  nand NAND2_4591(WX7705,II23582,II23583);
  nand NAND2_4592(II23588,WX7083,CRC_OUT_4_24);
  nand NAND2_4593(II23589,WX7083,II23588);
  nand NAND2_4594(II23590,CRC_OUT_4_24,II23588);
  nand NAND2_4595(WX7706,II23589,II23590);
  nand NAND2_4596(II23595,WX7084,CRC_OUT_4_23);
  nand NAND2_4597(II23596,WX7084,II23595);
  nand NAND2_4598(II23597,CRC_OUT_4_23,II23595);
  nand NAND2_4599(WX7707,II23596,II23597);
  nand NAND2_4600(II23602,WX7085,CRC_OUT_4_22);
  nand NAND2_4601(II23603,WX7085,II23602);
  nand NAND2_4602(II23604,CRC_OUT_4_22,II23602);
  nand NAND2_4603(WX7708,II23603,II23604);
  nand NAND2_4604(II23609,WX7086,CRC_OUT_4_21);
  nand NAND2_4605(II23610,WX7086,II23609);
  nand NAND2_4606(II23611,CRC_OUT_4_21,II23609);
  nand NAND2_4607(WX7709,II23610,II23611);
  nand NAND2_4608(II23616,WX7087,CRC_OUT_4_20);
  nand NAND2_4609(II23617,WX7087,II23616);
  nand NAND2_4610(II23618,CRC_OUT_4_20,II23616);
  nand NAND2_4611(WX7710,II23617,II23618);
  nand NAND2_4612(II23623,WX7088,CRC_OUT_4_19);
  nand NAND2_4613(II23624,WX7088,II23623);
  nand NAND2_4614(II23625,CRC_OUT_4_19,II23623);
  nand NAND2_4615(WX7711,II23624,II23625);
  nand NAND2_4616(II23630,WX7089,CRC_OUT_4_18);
  nand NAND2_4617(II23631,WX7089,II23630);
  nand NAND2_4618(II23632,CRC_OUT_4_18,II23630);
  nand NAND2_4619(WX7712,II23631,II23632);
  nand NAND2_4620(II23637,WX7090,CRC_OUT_4_17);
  nand NAND2_4621(II23638,WX7090,II23637);
  nand NAND2_4622(II23639,CRC_OUT_4_17,II23637);
  nand NAND2_4623(WX7713,II23638,II23639);
  nand NAND2_4624(II23644,WX7091,CRC_OUT_4_16);
  nand NAND2_4625(II23645,WX7091,II23644);
  nand NAND2_4626(II23646,CRC_OUT_4_16,II23644);
  nand NAND2_4627(WX7714,II23645,II23646);
  nand NAND2_4628(II23651,WX7093,CRC_OUT_4_14);
  nand NAND2_4629(II23652,WX7093,II23651);
  nand NAND2_4630(II23653,CRC_OUT_4_14,II23651);
  nand NAND2_4631(WX7715,II23652,II23653);
  nand NAND2_4632(II23658,WX7094,CRC_OUT_4_13);
  nand NAND2_4633(II23659,WX7094,II23658);
  nand NAND2_4634(II23660,CRC_OUT_4_13,II23658);
  nand NAND2_4635(WX7716,II23659,II23660);
  nand NAND2_4636(II23665,WX7095,CRC_OUT_4_12);
  nand NAND2_4637(II23666,WX7095,II23665);
  nand NAND2_4638(II23667,CRC_OUT_4_12,II23665);
  nand NAND2_4639(WX7717,II23666,II23667);
  nand NAND2_4640(II23672,WX7096,CRC_OUT_4_11);
  nand NAND2_4641(II23673,WX7096,II23672);
  nand NAND2_4642(II23674,CRC_OUT_4_11,II23672);
  nand NAND2_4643(WX7718,II23673,II23674);
  nand NAND2_4644(II23679,WX7098,CRC_OUT_4_9);
  nand NAND2_4645(II23680,WX7098,II23679);
  nand NAND2_4646(II23681,CRC_OUT_4_9,II23679);
  nand NAND2_4647(WX7719,II23680,II23681);
  nand NAND2_4648(II23686,WX7099,CRC_OUT_4_8);
  nand NAND2_4649(II23687,WX7099,II23686);
  nand NAND2_4650(II23688,CRC_OUT_4_8,II23686);
  nand NAND2_4651(WX7720,II23687,II23688);
  nand NAND2_4652(II23693,WX7100,CRC_OUT_4_7);
  nand NAND2_4653(II23694,WX7100,II23693);
  nand NAND2_4654(II23695,CRC_OUT_4_7,II23693);
  nand NAND2_4655(WX7721,II23694,II23695);
  nand NAND2_4656(II23700,WX7101,CRC_OUT_4_6);
  nand NAND2_4657(II23701,WX7101,II23700);
  nand NAND2_4658(II23702,CRC_OUT_4_6,II23700);
  nand NAND2_4659(WX7722,II23701,II23702);
  nand NAND2_4660(II23707,WX7102,CRC_OUT_4_5);
  nand NAND2_4661(II23708,WX7102,II23707);
  nand NAND2_4662(II23709,CRC_OUT_4_5,II23707);
  nand NAND2_4663(WX7723,II23708,II23709);
  nand NAND2_4664(II23714,WX7103,CRC_OUT_4_4);
  nand NAND2_4665(II23715,WX7103,II23714);
  nand NAND2_4666(II23716,CRC_OUT_4_4,II23714);
  nand NAND2_4667(WX7724,II23715,II23716);
  nand NAND2_4668(II23721,WX7105,CRC_OUT_4_2);
  nand NAND2_4669(II23722,WX7105,II23721);
  nand NAND2_4670(II23723,CRC_OUT_4_2,II23721);
  nand NAND2_4671(WX7725,II23722,II23723);
  nand NAND2_4672(II23728,WX7106,CRC_OUT_4_1);
  nand NAND2_4673(II23729,WX7106,II23728);
  nand NAND2_4674(II23730,CRC_OUT_4_1,II23728);
  nand NAND2_4675(WX7726,II23729,II23730);
  nand NAND2_4676(II23735,WX7107,CRC_OUT_4_0);
  nand NAND2_4677(II23736,WX7107,II23735);
  nand NAND2_4678(II23737,CRC_OUT_4_0,II23735);
  nand NAND2_4679(WX7727,II23736,II23737);
  nand NAND2_4680(II26018,WX8759,WX8403);
  nand NAND2_4681(II26019,WX8759,II26018);
  nand NAND2_4682(II26020,WX8403,II26018);
  nand NAND2_4683(II26017,II26019,II26020);
  nand NAND2_4684(II26025,WX8467,II26017);
  nand NAND2_4685(II26026,WX8467,II26025);
  nand NAND2_4686(II26027,II26017,II26025);
  nand NAND2_4687(II26016,II26026,II26027);
  nand NAND2_4688(II26033,WX8531,WX8595);
  nand NAND2_4689(II26034,WX8531,II26033);
  nand NAND2_4690(II26035,WX8595,II26033);
  nand NAND2_4691(II26032,II26034,II26035);
  nand NAND2_4692(II26040,II26016,II26032);
  nand NAND2_4693(II26041,II26016,II26040);
  nand NAND2_4694(II26042,II26032,II26040);
  nand NAND2_4695(WX8658,II26041,II26042);
  nand NAND2_4696(II26049,WX8759,WX8405);
  nand NAND2_4697(II26050,WX8759,II26049);
  nand NAND2_4698(II26051,WX8405,II26049);
  nand NAND2_4699(II26048,II26050,II26051);
  nand NAND2_4700(II26056,WX8469,II26048);
  nand NAND2_4701(II26057,WX8469,II26056);
  nand NAND2_4702(II26058,II26048,II26056);
  nand NAND2_4703(II26047,II26057,II26058);
  nand NAND2_4704(II26064,WX8533,WX8597);
  nand NAND2_4705(II26065,WX8533,II26064);
  nand NAND2_4706(II26066,WX8597,II26064);
  nand NAND2_4707(II26063,II26065,II26066);
  nand NAND2_4708(II26071,II26047,II26063);
  nand NAND2_4709(II26072,II26047,II26071);
  nand NAND2_4710(II26073,II26063,II26071);
  nand NAND2_4711(WX8659,II26072,II26073);
  nand NAND2_4712(II26080,WX8759,WX8407);
  nand NAND2_4713(II26081,WX8759,II26080);
  nand NAND2_4714(II26082,WX8407,II26080);
  nand NAND2_4715(II26079,II26081,II26082);
  nand NAND2_4716(II26087,WX8471,II26079);
  nand NAND2_4717(II26088,WX8471,II26087);
  nand NAND2_4718(II26089,II26079,II26087);
  nand NAND2_4719(II26078,II26088,II26089);
  nand NAND2_4720(II26095,WX8535,WX8599);
  nand NAND2_4721(II26096,WX8535,II26095);
  nand NAND2_4722(II26097,WX8599,II26095);
  nand NAND2_4723(II26094,II26096,II26097);
  nand NAND2_4724(II26102,II26078,II26094);
  nand NAND2_4725(II26103,II26078,II26102);
  nand NAND2_4726(II26104,II26094,II26102);
  nand NAND2_4727(WX8660,II26103,II26104);
  nand NAND2_4728(II26111,WX8759,WX8409);
  nand NAND2_4729(II26112,WX8759,II26111);
  nand NAND2_4730(II26113,WX8409,II26111);
  nand NAND2_4731(II26110,II26112,II26113);
  nand NAND2_4732(II26118,WX8473,II26110);
  nand NAND2_4733(II26119,WX8473,II26118);
  nand NAND2_4734(II26120,II26110,II26118);
  nand NAND2_4735(II26109,II26119,II26120);
  nand NAND2_4736(II26126,WX8537,WX8601);
  nand NAND2_4737(II26127,WX8537,II26126);
  nand NAND2_4738(II26128,WX8601,II26126);
  nand NAND2_4739(II26125,II26127,II26128);
  nand NAND2_4740(II26133,II26109,II26125);
  nand NAND2_4741(II26134,II26109,II26133);
  nand NAND2_4742(II26135,II26125,II26133);
  nand NAND2_4743(WX8661,II26134,II26135);
  nand NAND2_4744(II26142,WX8759,WX8411);
  nand NAND2_4745(II26143,WX8759,II26142);
  nand NAND2_4746(II26144,WX8411,II26142);
  nand NAND2_4747(II26141,II26143,II26144);
  nand NAND2_4748(II26149,WX8475,II26141);
  nand NAND2_4749(II26150,WX8475,II26149);
  nand NAND2_4750(II26151,II26141,II26149);
  nand NAND2_4751(II26140,II26150,II26151);
  nand NAND2_4752(II26157,WX8539,WX8603);
  nand NAND2_4753(II26158,WX8539,II26157);
  nand NAND2_4754(II26159,WX8603,II26157);
  nand NAND2_4755(II26156,II26158,II26159);
  nand NAND2_4756(II26164,II26140,II26156);
  nand NAND2_4757(II26165,II26140,II26164);
  nand NAND2_4758(II26166,II26156,II26164);
  nand NAND2_4759(WX8662,II26165,II26166);
  nand NAND2_4760(II26173,WX8759,WX8413);
  nand NAND2_4761(II26174,WX8759,II26173);
  nand NAND2_4762(II26175,WX8413,II26173);
  nand NAND2_4763(II26172,II26174,II26175);
  nand NAND2_4764(II26180,WX8477,II26172);
  nand NAND2_4765(II26181,WX8477,II26180);
  nand NAND2_4766(II26182,II26172,II26180);
  nand NAND2_4767(II26171,II26181,II26182);
  nand NAND2_4768(II26188,WX8541,WX8605);
  nand NAND2_4769(II26189,WX8541,II26188);
  nand NAND2_4770(II26190,WX8605,II26188);
  nand NAND2_4771(II26187,II26189,II26190);
  nand NAND2_4772(II26195,II26171,II26187);
  nand NAND2_4773(II26196,II26171,II26195);
  nand NAND2_4774(II26197,II26187,II26195);
  nand NAND2_4775(WX8663,II26196,II26197);
  nand NAND2_4776(II26204,WX8759,WX8415);
  nand NAND2_4777(II26205,WX8759,II26204);
  nand NAND2_4778(II26206,WX8415,II26204);
  nand NAND2_4779(II26203,II26205,II26206);
  nand NAND2_4780(II26211,WX8479,II26203);
  nand NAND2_4781(II26212,WX8479,II26211);
  nand NAND2_4782(II26213,II26203,II26211);
  nand NAND2_4783(II26202,II26212,II26213);
  nand NAND2_4784(II26219,WX8543,WX8607);
  nand NAND2_4785(II26220,WX8543,II26219);
  nand NAND2_4786(II26221,WX8607,II26219);
  nand NAND2_4787(II26218,II26220,II26221);
  nand NAND2_4788(II26226,II26202,II26218);
  nand NAND2_4789(II26227,II26202,II26226);
  nand NAND2_4790(II26228,II26218,II26226);
  nand NAND2_4791(WX8664,II26227,II26228);
  nand NAND2_4792(II26235,WX8759,WX8417);
  nand NAND2_4793(II26236,WX8759,II26235);
  nand NAND2_4794(II26237,WX8417,II26235);
  nand NAND2_4795(II26234,II26236,II26237);
  nand NAND2_4796(II26242,WX8481,II26234);
  nand NAND2_4797(II26243,WX8481,II26242);
  nand NAND2_4798(II26244,II26234,II26242);
  nand NAND2_4799(II26233,II26243,II26244);
  nand NAND2_4800(II26250,WX8545,WX8609);
  nand NAND2_4801(II26251,WX8545,II26250);
  nand NAND2_4802(II26252,WX8609,II26250);
  nand NAND2_4803(II26249,II26251,II26252);
  nand NAND2_4804(II26257,II26233,II26249);
  nand NAND2_4805(II26258,II26233,II26257);
  nand NAND2_4806(II26259,II26249,II26257);
  nand NAND2_4807(WX8665,II26258,II26259);
  nand NAND2_4808(II26266,WX8759,WX8419);
  nand NAND2_4809(II26267,WX8759,II26266);
  nand NAND2_4810(II26268,WX8419,II26266);
  nand NAND2_4811(II26265,II26267,II26268);
  nand NAND2_4812(II26273,WX8483,II26265);
  nand NAND2_4813(II26274,WX8483,II26273);
  nand NAND2_4814(II26275,II26265,II26273);
  nand NAND2_4815(II26264,II26274,II26275);
  nand NAND2_4816(II26281,WX8547,WX8611);
  nand NAND2_4817(II26282,WX8547,II26281);
  nand NAND2_4818(II26283,WX8611,II26281);
  nand NAND2_4819(II26280,II26282,II26283);
  nand NAND2_4820(II26288,II26264,II26280);
  nand NAND2_4821(II26289,II26264,II26288);
  nand NAND2_4822(II26290,II26280,II26288);
  nand NAND2_4823(WX8666,II26289,II26290);
  nand NAND2_4824(II26297,WX8759,WX8421);
  nand NAND2_4825(II26298,WX8759,II26297);
  nand NAND2_4826(II26299,WX8421,II26297);
  nand NAND2_4827(II26296,II26298,II26299);
  nand NAND2_4828(II26304,WX8485,II26296);
  nand NAND2_4829(II26305,WX8485,II26304);
  nand NAND2_4830(II26306,II26296,II26304);
  nand NAND2_4831(II26295,II26305,II26306);
  nand NAND2_4832(II26312,WX8549,WX8613);
  nand NAND2_4833(II26313,WX8549,II26312);
  nand NAND2_4834(II26314,WX8613,II26312);
  nand NAND2_4835(II26311,II26313,II26314);
  nand NAND2_4836(II26319,II26295,II26311);
  nand NAND2_4837(II26320,II26295,II26319);
  nand NAND2_4838(II26321,II26311,II26319);
  nand NAND2_4839(WX8667,II26320,II26321);
  nand NAND2_4840(II26328,WX8759,WX8423);
  nand NAND2_4841(II26329,WX8759,II26328);
  nand NAND2_4842(II26330,WX8423,II26328);
  nand NAND2_4843(II26327,II26329,II26330);
  nand NAND2_4844(II26335,WX8487,II26327);
  nand NAND2_4845(II26336,WX8487,II26335);
  nand NAND2_4846(II26337,II26327,II26335);
  nand NAND2_4847(II26326,II26336,II26337);
  nand NAND2_4848(II26343,WX8551,WX8615);
  nand NAND2_4849(II26344,WX8551,II26343);
  nand NAND2_4850(II26345,WX8615,II26343);
  nand NAND2_4851(II26342,II26344,II26345);
  nand NAND2_4852(II26350,II26326,II26342);
  nand NAND2_4853(II26351,II26326,II26350);
  nand NAND2_4854(II26352,II26342,II26350);
  nand NAND2_4855(WX8668,II26351,II26352);
  nand NAND2_4856(II26359,WX8759,WX8425);
  nand NAND2_4857(II26360,WX8759,II26359);
  nand NAND2_4858(II26361,WX8425,II26359);
  nand NAND2_4859(II26358,II26360,II26361);
  nand NAND2_4860(II26366,WX8489,II26358);
  nand NAND2_4861(II26367,WX8489,II26366);
  nand NAND2_4862(II26368,II26358,II26366);
  nand NAND2_4863(II26357,II26367,II26368);
  nand NAND2_4864(II26374,WX8553,WX8617);
  nand NAND2_4865(II26375,WX8553,II26374);
  nand NAND2_4866(II26376,WX8617,II26374);
  nand NAND2_4867(II26373,II26375,II26376);
  nand NAND2_4868(II26381,II26357,II26373);
  nand NAND2_4869(II26382,II26357,II26381);
  nand NAND2_4870(II26383,II26373,II26381);
  nand NAND2_4871(WX8669,II26382,II26383);
  nand NAND2_4872(II26390,WX8759,WX8427);
  nand NAND2_4873(II26391,WX8759,II26390);
  nand NAND2_4874(II26392,WX8427,II26390);
  nand NAND2_4875(II26389,II26391,II26392);
  nand NAND2_4876(II26397,WX8491,II26389);
  nand NAND2_4877(II26398,WX8491,II26397);
  nand NAND2_4878(II26399,II26389,II26397);
  nand NAND2_4879(II26388,II26398,II26399);
  nand NAND2_4880(II26405,WX8555,WX8619);
  nand NAND2_4881(II26406,WX8555,II26405);
  nand NAND2_4882(II26407,WX8619,II26405);
  nand NAND2_4883(II26404,II26406,II26407);
  nand NAND2_4884(II26412,II26388,II26404);
  nand NAND2_4885(II26413,II26388,II26412);
  nand NAND2_4886(II26414,II26404,II26412);
  nand NAND2_4887(WX8670,II26413,II26414);
  nand NAND2_4888(II26421,WX8759,WX8429);
  nand NAND2_4889(II26422,WX8759,II26421);
  nand NAND2_4890(II26423,WX8429,II26421);
  nand NAND2_4891(II26420,II26422,II26423);
  nand NAND2_4892(II26428,WX8493,II26420);
  nand NAND2_4893(II26429,WX8493,II26428);
  nand NAND2_4894(II26430,II26420,II26428);
  nand NAND2_4895(II26419,II26429,II26430);
  nand NAND2_4896(II26436,WX8557,WX8621);
  nand NAND2_4897(II26437,WX8557,II26436);
  nand NAND2_4898(II26438,WX8621,II26436);
  nand NAND2_4899(II26435,II26437,II26438);
  nand NAND2_4900(II26443,II26419,II26435);
  nand NAND2_4901(II26444,II26419,II26443);
  nand NAND2_4902(II26445,II26435,II26443);
  nand NAND2_4903(WX8671,II26444,II26445);
  nand NAND2_4904(II26452,WX8759,WX8431);
  nand NAND2_4905(II26453,WX8759,II26452);
  nand NAND2_4906(II26454,WX8431,II26452);
  nand NAND2_4907(II26451,II26453,II26454);
  nand NAND2_4908(II26459,WX8495,II26451);
  nand NAND2_4909(II26460,WX8495,II26459);
  nand NAND2_4910(II26461,II26451,II26459);
  nand NAND2_4911(II26450,II26460,II26461);
  nand NAND2_4912(II26467,WX8559,WX8623);
  nand NAND2_4913(II26468,WX8559,II26467);
  nand NAND2_4914(II26469,WX8623,II26467);
  nand NAND2_4915(II26466,II26468,II26469);
  nand NAND2_4916(II26474,II26450,II26466);
  nand NAND2_4917(II26475,II26450,II26474);
  nand NAND2_4918(II26476,II26466,II26474);
  nand NAND2_4919(WX8672,II26475,II26476);
  nand NAND2_4920(II26483,WX8759,WX8433);
  nand NAND2_4921(II26484,WX8759,II26483);
  nand NAND2_4922(II26485,WX8433,II26483);
  nand NAND2_4923(II26482,II26484,II26485);
  nand NAND2_4924(II26490,WX8497,II26482);
  nand NAND2_4925(II26491,WX8497,II26490);
  nand NAND2_4926(II26492,II26482,II26490);
  nand NAND2_4927(II26481,II26491,II26492);
  nand NAND2_4928(II26498,WX8561,WX8625);
  nand NAND2_4929(II26499,WX8561,II26498);
  nand NAND2_4930(II26500,WX8625,II26498);
  nand NAND2_4931(II26497,II26499,II26500);
  nand NAND2_4932(II26505,II26481,II26497);
  nand NAND2_4933(II26506,II26481,II26505);
  nand NAND2_4934(II26507,II26497,II26505);
  nand NAND2_4935(WX8673,II26506,II26507);
  nand NAND2_4936(II26514,WX8760,WX8435);
  nand NAND2_4937(II26515,WX8760,II26514);
  nand NAND2_4938(II26516,WX8435,II26514);
  nand NAND2_4939(II26513,II26515,II26516);
  nand NAND2_4940(II26521,WX8499,II26513);
  nand NAND2_4941(II26522,WX8499,II26521);
  nand NAND2_4942(II26523,II26513,II26521);
  nand NAND2_4943(II26512,II26522,II26523);
  nand NAND2_4944(II26529,WX8563,WX8627);
  nand NAND2_4945(II26530,WX8563,II26529);
  nand NAND2_4946(II26531,WX8627,II26529);
  nand NAND2_4947(II26528,II26530,II26531);
  nand NAND2_4948(II26536,II26512,II26528);
  nand NAND2_4949(II26537,II26512,II26536);
  nand NAND2_4950(II26538,II26528,II26536);
  nand NAND2_4951(WX8674,II26537,II26538);
  nand NAND2_4952(II26545,WX8760,WX8437);
  nand NAND2_4953(II26546,WX8760,II26545);
  nand NAND2_4954(II26547,WX8437,II26545);
  nand NAND2_4955(II26544,II26546,II26547);
  nand NAND2_4956(II26552,WX8501,II26544);
  nand NAND2_4957(II26553,WX8501,II26552);
  nand NAND2_4958(II26554,II26544,II26552);
  nand NAND2_4959(II26543,II26553,II26554);
  nand NAND2_4960(II26560,WX8565,WX8629);
  nand NAND2_4961(II26561,WX8565,II26560);
  nand NAND2_4962(II26562,WX8629,II26560);
  nand NAND2_4963(II26559,II26561,II26562);
  nand NAND2_4964(II26567,II26543,II26559);
  nand NAND2_4965(II26568,II26543,II26567);
  nand NAND2_4966(II26569,II26559,II26567);
  nand NAND2_4967(WX8675,II26568,II26569);
  nand NAND2_4968(II26576,WX8760,WX8439);
  nand NAND2_4969(II26577,WX8760,II26576);
  nand NAND2_4970(II26578,WX8439,II26576);
  nand NAND2_4971(II26575,II26577,II26578);
  nand NAND2_4972(II26583,WX8503,II26575);
  nand NAND2_4973(II26584,WX8503,II26583);
  nand NAND2_4974(II26585,II26575,II26583);
  nand NAND2_4975(II26574,II26584,II26585);
  nand NAND2_4976(II26591,WX8567,WX8631);
  nand NAND2_4977(II26592,WX8567,II26591);
  nand NAND2_4978(II26593,WX8631,II26591);
  nand NAND2_4979(II26590,II26592,II26593);
  nand NAND2_4980(II26598,II26574,II26590);
  nand NAND2_4981(II26599,II26574,II26598);
  nand NAND2_4982(II26600,II26590,II26598);
  nand NAND2_4983(WX8676,II26599,II26600);
  nand NAND2_4984(II26607,WX8760,WX8441);
  nand NAND2_4985(II26608,WX8760,II26607);
  nand NAND2_4986(II26609,WX8441,II26607);
  nand NAND2_4987(II26606,II26608,II26609);
  nand NAND2_4988(II26614,WX8505,II26606);
  nand NAND2_4989(II26615,WX8505,II26614);
  nand NAND2_4990(II26616,II26606,II26614);
  nand NAND2_4991(II26605,II26615,II26616);
  nand NAND2_4992(II26622,WX8569,WX8633);
  nand NAND2_4993(II26623,WX8569,II26622);
  nand NAND2_4994(II26624,WX8633,II26622);
  nand NAND2_4995(II26621,II26623,II26624);
  nand NAND2_4996(II26629,II26605,II26621);
  nand NAND2_4997(II26630,II26605,II26629);
  nand NAND2_4998(II26631,II26621,II26629);
  nand NAND2_4999(WX8677,II26630,II26631);
  nand NAND2_5000(II26638,WX8760,WX8443);
  nand NAND2_5001(II26639,WX8760,II26638);
  nand NAND2_5002(II26640,WX8443,II26638);
  nand NAND2_5003(II26637,II26639,II26640);
  nand NAND2_5004(II26645,WX8507,II26637);
  nand NAND2_5005(II26646,WX8507,II26645);
  nand NAND2_5006(II26647,II26637,II26645);
  nand NAND2_5007(II26636,II26646,II26647);
  nand NAND2_5008(II26653,WX8571,WX8635);
  nand NAND2_5009(II26654,WX8571,II26653);
  nand NAND2_5010(II26655,WX8635,II26653);
  nand NAND2_5011(II26652,II26654,II26655);
  nand NAND2_5012(II26660,II26636,II26652);
  nand NAND2_5013(II26661,II26636,II26660);
  nand NAND2_5014(II26662,II26652,II26660);
  nand NAND2_5015(WX8678,II26661,II26662);
  nand NAND2_5016(II26669,WX8760,WX8445);
  nand NAND2_5017(II26670,WX8760,II26669);
  nand NAND2_5018(II26671,WX8445,II26669);
  nand NAND2_5019(II26668,II26670,II26671);
  nand NAND2_5020(II26676,WX8509,II26668);
  nand NAND2_5021(II26677,WX8509,II26676);
  nand NAND2_5022(II26678,II26668,II26676);
  nand NAND2_5023(II26667,II26677,II26678);
  nand NAND2_5024(II26684,WX8573,WX8637);
  nand NAND2_5025(II26685,WX8573,II26684);
  nand NAND2_5026(II26686,WX8637,II26684);
  nand NAND2_5027(II26683,II26685,II26686);
  nand NAND2_5028(II26691,II26667,II26683);
  nand NAND2_5029(II26692,II26667,II26691);
  nand NAND2_5030(II26693,II26683,II26691);
  nand NAND2_5031(WX8679,II26692,II26693);
  nand NAND2_5032(II26700,WX8760,WX8447);
  nand NAND2_5033(II26701,WX8760,II26700);
  nand NAND2_5034(II26702,WX8447,II26700);
  nand NAND2_5035(II26699,II26701,II26702);
  nand NAND2_5036(II26707,WX8511,II26699);
  nand NAND2_5037(II26708,WX8511,II26707);
  nand NAND2_5038(II26709,II26699,II26707);
  nand NAND2_5039(II26698,II26708,II26709);
  nand NAND2_5040(II26715,WX8575,WX8639);
  nand NAND2_5041(II26716,WX8575,II26715);
  nand NAND2_5042(II26717,WX8639,II26715);
  nand NAND2_5043(II26714,II26716,II26717);
  nand NAND2_5044(II26722,II26698,II26714);
  nand NAND2_5045(II26723,II26698,II26722);
  nand NAND2_5046(II26724,II26714,II26722);
  nand NAND2_5047(WX8680,II26723,II26724);
  nand NAND2_5048(II26731,WX8760,WX8449);
  nand NAND2_5049(II26732,WX8760,II26731);
  nand NAND2_5050(II26733,WX8449,II26731);
  nand NAND2_5051(II26730,II26732,II26733);
  nand NAND2_5052(II26738,WX8513,II26730);
  nand NAND2_5053(II26739,WX8513,II26738);
  nand NAND2_5054(II26740,II26730,II26738);
  nand NAND2_5055(II26729,II26739,II26740);
  nand NAND2_5056(II26746,WX8577,WX8641);
  nand NAND2_5057(II26747,WX8577,II26746);
  nand NAND2_5058(II26748,WX8641,II26746);
  nand NAND2_5059(II26745,II26747,II26748);
  nand NAND2_5060(II26753,II26729,II26745);
  nand NAND2_5061(II26754,II26729,II26753);
  nand NAND2_5062(II26755,II26745,II26753);
  nand NAND2_5063(WX8681,II26754,II26755);
  nand NAND2_5064(II26762,WX8760,WX8451);
  nand NAND2_5065(II26763,WX8760,II26762);
  nand NAND2_5066(II26764,WX8451,II26762);
  nand NAND2_5067(II26761,II26763,II26764);
  nand NAND2_5068(II26769,WX8515,II26761);
  nand NAND2_5069(II26770,WX8515,II26769);
  nand NAND2_5070(II26771,II26761,II26769);
  nand NAND2_5071(II26760,II26770,II26771);
  nand NAND2_5072(II26777,WX8579,WX8643);
  nand NAND2_5073(II26778,WX8579,II26777);
  nand NAND2_5074(II26779,WX8643,II26777);
  nand NAND2_5075(II26776,II26778,II26779);
  nand NAND2_5076(II26784,II26760,II26776);
  nand NAND2_5077(II26785,II26760,II26784);
  nand NAND2_5078(II26786,II26776,II26784);
  nand NAND2_5079(WX8682,II26785,II26786);
  nand NAND2_5080(II26793,WX8760,WX8453);
  nand NAND2_5081(II26794,WX8760,II26793);
  nand NAND2_5082(II26795,WX8453,II26793);
  nand NAND2_5083(II26792,II26794,II26795);
  nand NAND2_5084(II26800,WX8517,II26792);
  nand NAND2_5085(II26801,WX8517,II26800);
  nand NAND2_5086(II26802,II26792,II26800);
  nand NAND2_5087(II26791,II26801,II26802);
  nand NAND2_5088(II26808,WX8581,WX8645);
  nand NAND2_5089(II26809,WX8581,II26808);
  nand NAND2_5090(II26810,WX8645,II26808);
  nand NAND2_5091(II26807,II26809,II26810);
  nand NAND2_5092(II26815,II26791,II26807);
  nand NAND2_5093(II26816,II26791,II26815);
  nand NAND2_5094(II26817,II26807,II26815);
  nand NAND2_5095(WX8683,II26816,II26817);
  nand NAND2_5096(II26824,WX8760,WX8455);
  nand NAND2_5097(II26825,WX8760,II26824);
  nand NAND2_5098(II26826,WX8455,II26824);
  nand NAND2_5099(II26823,II26825,II26826);
  nand NAND2_5100(II26831,WX8519,II26823);
  nand NAND2_5101(II26832,WX8519,II26831);
  nand NAND2_5102(II26833,II26823,II26831);
  nand NAND2_5103(II26822,II26832,II26833);
  nand NAND2_5104(II26839,WX8583,WX8647);
  nand NAND2_5105(II26840,WX8583,II26839);
  nand NAND2_5106(II26841,WX8647,II26839);
  nand NAND2_5107(II26838,II26840,II26841);
  nand NAND2_5108(II26846,II26822,II26838);
  nand NAND2_5109(II26847,II26822,II26846);
  nand NAND2_5110(II26848,II26838,II26846);
  nand NAND2_5111(WX8684,II26847,II26848);
  nand NAND2_5112(II26855,WX8760,WX8457);
  nand NAND2_5113(II26856,WX8760,II26855);
  nand NAND2_5114(II26857,WX8457,II26855);
  nand NAND2_5115(II26854,II26856,II26857);
  nand NAND2_5116(II26862,WX8521,II26854);
  nand NAND2_5117(II26863,WX8521,II26862);
  nand NAND2_5118(II26864,II26854,II26862);
  nand NAND2_5119(II26853,II26863,II26864);
  nand NAND2_5120(II26870,WX8585,WX8649);
  nand NAND2_5121(II26871,WX8585,II26870);
  nand NAND2_5122(II26872,WX8649,II26870);
  nand NAND2_5123(II26869,II26871,II26872);
  nand NAND2_5124(II26877,II26853,II26869);
  nand NAND2_5125(II26878,II26853,II26877);
  nand NAND2_5126(II26879,II26869,II26877);
  nand NAND2_5127(WX8685,II26878,II26879);
  nand NAND2_5128(II26886,WX8760,WX8459);
  nand NAND2_5129(II26887,WX8760,II26886);
  nand NAND2_5130(II26888,WX8459,II26886);
  nand NAND2_5131(II26885,II26887,II26888);
  nand NAND2_5132(II26893,WX8523,II26885);
  nand NAND2_5133(II26894,WX8523,II26893);
  nand NAND2_5134(II26895,II26885,II26893);
  nand NAND2_5135(II26884,II26894,II26895);
  nand NAND2_5136(II26901,WX8587,WX8651);
  nand NAND2_5137(II26902,WX8587,II26901);
  nand NAND2_5138(II26903,WX8651,II26901);
  nand NAND2_5139(II26900,II26902,II26903);
  nand NAND2_5140(II26908,II26884,II26900);
  nand NAND2_5141(II26909,II26884,II26908);
  nand NAND2_5142(II26910,II26900,II26908);
  nand NAND2_5143(WX8686,II26909,II26910);
  nand NAND2_5144(II26917,WX8760,WX8461);
  nand NAND2_5145(II26918,WX8760,II26917);
  nand NAND2_5146(II26919,WX8461,II26917);
  nand NAND2_5147(II26916,II26918,II26919);
  nand NAND2_5148(II26924,WX8525,II26916);
  nand NAND2_5149(II26925,WX8525,II26924);
  nand NAND2_5150(II26926,II26916,II26924);
  nand NAND2_5151(II26915,II26925,II26926);
  nand NAND2_5152(II26932,WX8589,WX8653);
  nand NAND2_5153(II26933,WX8589,II26932);
  nand NAND2_5154(II26934,WX8653,II26932);
  nand NAND2_5155(II26931,II26933,II26934);
  nand NAND2_5156(II26939,II26915,II26931);
  nand NAND2_5157(II26940,II26915,II26939);
  nand NAND2_5158(II26941,II26931,II26939);
  nand NAND2_5159(WX8687,II26940,II26941);
  nand NAND2_5160(II26948,WX8760,WX8463);
  nand NAND2_5161(II26949,WX8760,II26948);
  nand NAND2_5162(II26950,WX8463,II26948);
  nand NAND2_5163(II26947,II26949,II26950);
  nand NAND2_5164(II26955,WX8527,II26947);
  nand NAND2_5165(II26956,WX8527,II26955);
  nand NAND2_5166(II26957,II26947,II26955);
  nand NAND2_5167(II26946,II26956,II26957);
  nand NAND2_5168(II26963,WX8591,WX8655);
  nand NAND2_5169(II26964,WX8591,II26963);
  nand NAND2_5170(II26965,WX8655,II26963);
  nand NAND2_5171(II26962,II26964,II26965);
  nand NAND2_5172(II26970,II26946,II26962);
  nand NAND2_5173(II26971,II26946,II26970);
  nand NAND2_5174(II26972,II26962,II26970);
  nand NAND2_5175(WX8688,II26971,II26972);
  nand NAND2_5176(II26979,WX8760,WX8465);
  nand NAND2_5177(II26980,WX8760,II26979);
  nand NAND2_5178(II26981,WX8465,II26979);
  nand NAND2_5179(II26978,II26980,II26981);
  nand NAND2_5180(II26986,WX8529,II26978);
  nand NAND2_5181(II26987,WX8529,II26986);
  nand NAND2_5182(II26988,II26978,II26986);
  nand NAND2_5183(II26977,II26987,II26988);
  nand NAND2_5184(II26994,WX8593,WX8657);
  nand NAND2_5185(II26995,WX8593,II26994);
  nand NAND2_5186(II26996,WX8657,II26994);
  nand NAND2_5187(II26993,II26995,II26996);
  nand NAND2_5188(II27001,II26977,II26993);
  nand NAND2_5189(II27002,II26977,II27001);
  nand NAND2_5190(II27003,II26993,II27001);
  nand NAND2_5191(WX8689,II27002,II27003);
  nand NAND2_5192(II27082,WX8338,WX8243);
  nand NAND2_5193(II27083,WX8338,II27082);
  nand NAND2_5194(II27084,WX8243,II27082);
  nand NAND2_5195(WX8764,II27083,II27084);
  nand NAND2_5196(II27095,WX8339,WX8245);
  nand NAND2_5197(II27096,WX8339,II27095);
  nand NAND2_5198(II27097,WX8245,II27095);
  nand NAND2_5199(WX8771,II27096,II27097);
  nand NAND2_5200(II27108,WX8340,WX8247);
  nand NAND2_5201(II27109,WX8340,II27108);
  nand NAND2_5202(II27110,WX8247,II27108);
  nand NAND2_5203(WX8778,II27109,II27110);
  nand NAND2_5204(II27121,WX8341,WX8249);
  nand NAND2_5205(II27122,WX8341,II27121);
  nand NAND2_5206(II27123,WX8249,II27121);
  nand NAND2_5207(WX8785,II27122,II27123);
  nand NAND2_5208(II27134,WX8342,WX8251);
  nand NAND2_5209(II27135,WX8342,II27134);
  nand NAND2_5210(II27136,WX8251,II27134);
  nand NAND2_5211(WX8792,II27135,II27136);
  nand NAND2_5212(II27147,WX8343,WX8253);
  nand NAND2_5213(II27148,WX8343,II27147);
  nand NAND2_5214(II27149,WX8253,II27147);
  nand NAND2_5215(WX8799,II27148,II27149);
  nand NAND2_5216(II27160,WX8344,WX8255);
  nand NAND2_5217(II27161,WX8344,II27160);
  nand NAND2_5218(II27162,WX8255,II27160);
  nand NAND2_5219(WX8806,II27161,II27162);
  nand NAND2_5220(II27173,WX8345,WX8257);
  nand NAND2_5221(II27174,WX8345,II27173);
  nand NAND2_5222(II27175,WX8257,II27173);
  nand NAND2_5223(WX8813,II27174,II27175);
  nand NAND2_5224(II27186,WX8346,WX8259);
  nand NAND2_5225(II27187,WX8346,II27186);
  nand NAND2_5226(II27188,WX8259,II27186);
  nand NAND2_5227(WX8820,II27187,II27188);
  nand NAND2_5228(II27199,WX8347,WX8261);
  nand NAND2_5229(II27200,WX8347,II27199);
  nand NAND2_5230(II27201,WX8261,II27199);
  nand NAND2_5231(WX8827,II27200,II27201);
  nand NAND2_5232(II27212,WX8348,WX8263);
  nand NAND2_5233(II27213,WX8348,II27212);
  nand NAND2_5234(II27214,WX8263,II27212);
  nand NAND2_5235(WX8834,II27213,II27214);
  nand NAND2_5236(II27225,WX8349,WX8265);
  nand NAND2_5237(II27226,WX8349,II27225);
  nand NAND2_5238(II27227,WX8265,II27225);
  nand NAND2_5239(WX8841,II27226,II27227);
  nand NAND2_5240(II27238,WX8350,WX8267);
  nand NAND2_5241(II27239,WX8350,II27238);
  nand NAND2_5242(II27240,WX8267,II27238);
  nand NAND2_5243(WX8848,II27239,II27240);
  nand NAND2_5244(II27251,WX8351,WX8269);
  nand NAND2_5245(II27252,WX8351,II27251);
  nand NAND2_5246(II27253,WX8269,II27251);
  nand NAND2_5247(WX8855,II27252,II27253);
  nand NAND2_5248(II27264,WX8352,WX8271);
  nand NAND2_5249(II27265,WX8352,II27264);
  nand NAND2_5250(II27266,WX8271,II27264);
  nand NAND2_5251(WX8862,II27265,II27266);
  nand NAND2_5252(II27277,WX8353,WX8273);
  nand NAND2_5253(II27278,WX8353,II27277);
  nand NAND2_5254(II27279,WX8273,II27277);
  nand NAND2_5255(WX8869,II27278,II27279);
  nand NAND2_5256(II27290,WX8354,WX8275);
  nand NAND2_5257(II27291,WX8354,II27290);
  nand NAND2_5258(II27292,WX8275,II27290);
  nand NAND2_5259(WX8876,II27291,II27292);
  nand NAND2_5260(II27303,WX8355,WX8277);
  nand NAND2_5261(II27304,WX8355,II27303);
  nand NAND2_5262(II27305,WX8277,II27303);
  nand NAND2_5263(WX8883,II27304,II27305);
  nand NAND2_5264(II27316,WX8356,WX8279);
  nand NAND2_5265(II27317,WX8356,II27316);
  nand NAND2_5266(II27318,WX8279,II27316);
  nand NAND2_5267(WX8890,II27317,II27318);
  nand NAND2_5268(II27329,WX8357,WX8281);
  nand NAND2_5269(II27330,WX8357,II27329);
  nand NAND2_5270(II27331,WX8281,II27329);
  nand NAND2_5271(WX8897,II27330,II27331);
  nand NAND2_5272(II27342,WX8358,WX8283);
  nand NAND2_5273(II27343,WX8358,II27342);
  nand NAND2_5274(II27344,WX8283,II27342);
  nand NAND2_5275(WX8904,II27343,II27344);
  nand NAND2_5276(II27355,WX8359,WX8285);
  nand NAND2_5277(II27356,WX8359,II27355);
  nand NAND2_5278(II27357,WX8285,II27355);
  nand NAND2_5279(WX8911,II27356,II27357);
  nand NAND2_5280(II27368,WX8360,WX8287);
  nand NAND2_5281(II27369,WX8360,II27368);
  nand NAND2_5282(II27370,WX8287,II27368);
  nand NAND2_5283(WX8918,II27369,II27370);
  nand NAND2_5284(II27381,WX8361,WX8289);
  nand NAND2_5285(II27382,WX8361,II27381);
  nand NAND2_5286(II27383,WX8289,II27381);
  nand NAND2_5287(WX8925,II27382,II27383);
  nand NAND2_5288(II27394,WX8362,WX8291);
  nand NAND2_5289(II27395,WX8362,II27394);
  nand NAND2_5290(II27396,WX8291,II27394);
  nand NAND2_5291(WX8932,II27395,II27396);
  nand NAND2_5292(II27407,WX8363,WX8293);
  nand NAND2_5293(II27408,WX8363,II27407);
  nand NAND2_5294(II27409,WX8293,II27407);
  nand NAND2_5295(WX8939,II27408,II27409);
  nand NAND2_5296(II27420,WX8364,WX8295);
  nand NAND2_5297(II27421,WX8364,II27420);
  nand NAND2_5298(II27422,WX8295,II27420);
  nand NAND2_5299(WX8946,II27421,II27422);
  nand NAND2_5300(II27433,WX8365,WX8297);
  nand NAND2_5301(II27434,WX8365,II27433);
  nand NAND2_5302(II27435,WX8297,II27433);
  nand NAND2_5303(WX8953,II27434,II27435);
  nand NAND2_5304(II27446,WX8366,WX8299);
  nand NAND2_5305(II27447,WX8366,II27446);
  nand NAND2_5306(II27448,WX8299,II27446);
  nand NAND2_5307(WX8960,II27447,II27448);
  nand NAND2_5308(II27459,WX8367,WX8301);
  nand NAND2_5309(II27460,WX8367,II27459);
  nand NAND2_5310(II27461,WX8301,II27459);
  nand NAND2_5311(WX8967,II27460,II27461);
  nand NAND2_5312(II27472,WX8368,WX8303);
  nand NAND2_5313(II27473,WX8368,II27472);
  nand NAND2_5314(II27474,WX8303,II27472);
  nand NAND2_5315(WX8974,II27473,II27474);
  nand NAND2_5316(II27485,WX8369,WX8305);
  nand NAND2_5317(II27486,WX8369,II27485);
  nand NAND2_5318(II27487,WX8305,II27485);
  nand NAND2_5319(WX8981,II27486,II27487);
  nand NAND2_5320(II27500,WX8385,CRC_OUT_3_31);
  nand NAND2_5321(II27501,WX8385,II27500);
  nand NAND2_5322(II27502,CRC_OUT_3_31,II27500);
  nand NAND2_5323(II27499,II27501,II27502);
  nand NAND2_5324(II27507,CRC_OUT_3_15,II27499);
  nand NAND2_5325(II27508,CRC_OUT_3_15,II27507);
  nand NAND2_5326(II27509,II27499,II27507);
  nand NAND2_5327(WX8989,II27508,II27509);
  nand NAND2_5328(II27515,WX8390,CRC_OUT_3_31);
  nand NAND2_5329(II27516,WX8390,II27515);
  nand NAND2_5330(II27517,CRC_OUT_3_31,II27515);
  nand NAND2_5331(II27514,II27516,II27517);
  nand NAND2_5332(II27522,CRC_OUT_3_10,II27514);
  nand NAND2_5333(II27523,CRC_OUT_3_10,II27522);
  nand NAND2_5334(II27524,II27514,II27522);
  nand NAND2_5335(WX8990,II27523,II27524);
  nand NAND2_5336(II27530,WX8397,CRC_OUT_3_31);
  nand NAND2_5337(II27531,WX8397,II27530);
  nand NAND2_5338(II27532,CRC_OUT_3_31,II27530);
  nand NAND2_5339(II27529,II27531,II27532);
  nand NAND2_5340(II27537,CRC_OUT_3_3,II27529);
  nand NAND2_5341(II27538,CRC_OUT_3_3,II27537);
  nand NAND2_5342(II27539,II27529,II27537);
  nand NAND2_5343(WX8991,II27538,II27539);
  nand NAND2_5344(II27544,WX8401,CRC_OUT_3_31);
  nand NAND2_5345(II27545,WX8401,II27544);
  nand NAND2_5346(II27546,CRC_OUT_3_31,II27544);
  nand NAND2_5347(WX8992,II27545,II27546);
  nand NAND2_5348(II27551,WX8370,CRC_OUT_3_30);
  nand NAND2_5349(II27552,WX8370,II27551);
  nand NAND2_5350(II27553,CRC_OUT_3_30,II27551);
  nand NAND2_5351(WX8993,II27552,II27553);
  nand NAND2_5352(II27558,WX8371,CRC_OUT_3_29);
  nand NAND2_5353(II27559,WX8371,II27558);
  nand NAND2_5354(II27560,CRC_OUT_3_29,II27558);
  nand NAND2_5355(WX8994,II27559,II27560);
  nand NAND2_5356(II27565,WX8372,CRC_OUT_3_28);
  nand NAND2_5357(II27566,WX8372,II27565);
  nand NAND2_5358(II27567,CRC_OUT_3_28,II27565);
  nand NAND2_5359(WX8995,II27566,II27567);
  nand NAND2_5360(II27572,WX8373,CRC_OUT_3_27);
  nand NAND2_5361(II27573,WX8373,II27572);
  nand NAND2_5362(II27574,CRC_OUT_3_27,II27572);
  nand NAND2_5363(WX8996,II27573,II27574);
  nand NAND2_5364(II27579,WX8374,CRC_OUT_3_26);
  nand NAND2_5365(II27580,WX8374,II27579);
  nand NAND2_5366(II27581,CRC_OUT_3_26,II27579);
  nand NAND2_5367(WX8997,II27580,II27581);
  nand NAND2_5368(II27586,WX8375,CRC_OUT_3_25);
  nand NAND2_5369(II27587,WX8375,II27586);
  nand NAND2_5370(II27588,CRC_OUT_3_25,II27586);
  nand NAND2_5371(WX8998,II27587,II27588);
  nand NAND2_5372(II27593,WX8376,CRC_OUT_3_24);
  nand NAND2_5373(II27594,WX8376,II27593);
  nand NAND2_5374(II27595,CRC_OUT_3_24,II27593);
  nand NAND2_5375(WX8999,II27594,II27595);
  nand NAND2_5376(II27600,WX8377,CRC_OUT_3_23);
  nand NAND2_5377(II27601,WX8377,II27600);
  nand NAND2_5378(II27602,CRC_OUT_3_23,II27600);
  nand NAND2_5379(WX9000,II27601,II27602);
  nand NAND2_5380(II27607,WX8378,CRC_OUT_3_22);
  nand NAND2_5381(II27608,WX8378,II27607);
  nand NAND2_5382(II27609,CRC_OUT_3_22,II27607);
  nand NAND2_5383(WX9001,II27608,II27609);
  nand NAND2_5384(II27614,WX8379,CRC_OUT_3_21);
  nand NAND2_5385(II27615,WX8379,II27614);
  nand NAND2_5386(II27616,CRC_OUT_3_21,II27614);
  nand NAND2_5387(WX9002,II27615,II27616);
  nand NAND2_5388(II27621,WX8380,CRC_OUT_3_20);
  nand NAND2_5389(II27622,WX8380,II27621);
  nand NAND2_5390(II27623,CRC_OUT_3_20,II27621);
  nand NAND2_5391(WX9003,II27622,II27623);
  nand NAND2_5392(II27628,WX8381,CRC_OUT_3_19);
  nand NAND2_5393(II27629,WX8381,II27628);
  nand NAND2_5394(II27630,CRC_OUT_3_19,II27628);
  nand NAND2_5395(WX9004,II27629,II27630);
  nand NAND2_5396(II27635,WX8382,CRC_OUT_3_18);
  nand NAND2_5397(II27636,WX8382,II27635);
  nand NAND2_5398(II27637,CRC_OUT_3_18,II27635);
  nand NAND2_5399(WX9005,II27636,II27637);
  nand NAND2_5400(II27642,WX8383,CRC_OUT_3_17);
  nand NAND2_5401(II27643,WX8383,II27642);
  nand NAND2_5402(II27644,CRC_OUT_3_17,II27642);
  nand NAND2_5403(WX9006,II27643,II27644);
  nand NAND2_5404(II27649,WX8384,CRC_OUT_3_16);
  nand NAND2_5405(II27650,WX8384,II27649);
  nand NAND2_5406(II27651,CRC_OUT_3_16,II27649);
  nand NAND2_5407(WX9007,II27650,II27651);
  nand NAND2_5408(II27656,WX8386,CRC_OUT_3_14);
  nand NAND2_5409(II27657,WX8386,II27656);
  nand NAND2_5410(II27658,CRC_OUT_3_14,II27656);
  nand NAND2_5411(WX9008,II27657,II27658);
  nand NAND2_5412(II27663,WX8387,CRC_OUT_3_13);
  nand NAND2_5413(II27664,WX8387,II27663);
  nand NAND2_5414(II27665,CRC_OUT_3_13,II27663);
  nand NAND2_5415(WX9009,II27664,II27665);
  nand NAND2_5416(II27670,WX8388,CRC_OUT_3_12);
  nand NAND2_5417(II27671,WX8388,II27670);
  nand NAND2_5418(II27672,CRC_OUT_3_12,II27670);
  nand NAND2_5419(WX9010,II27671,II27672);
  nand NAND2_5420(II27677,WX8389,CRC_OUT_3_11);
  nand NAND2_5421(II27678,WX8389,II27677);
  nand NAND2_5422(II27679,CRC_OUT_3_11,II27677);
  nand NAND2_5423(WX9011,II27678,II27679);
  nand NAND2_5424(II27684,WX8391,CRC_OUT_3_9);
  nand NAND2_5425(II27685,WX8391,II27684);
  nand NAND2_5426(II27686,CRC_OUT_3_9,II27684);
  nand NAND2_5427(WX9012,II27685,II27686);
  nand NAND2_5428(II27691,WX8392,CRC_OUT_3_8);
  nand NAND2_5429(II27692,WX8392,II27691);
  nand NAND2_5430(II27693,CRC_OUT_3_8,II27691);
  nand NAND2_5431(WX9013,II27692,II27693);
  nand NAND2_5432(II27698,WX8393,CRC_OUT_3_7);
  nand NAND2_5433(II27699,WX8393,II27698);
  nand NAND2_5434(II27700,CRC_OUT_3_7,II27698);
  nand NAND2_5435(WX9014,II27699,II27700);
  nand NAND2_5436(II27705,WX8394,CRC_OUT_3_6);
  nand NAND2_5437(II27706,WX8394,II27705);
  nand NAND2_5438(II27707,CRC_OUT_3_6,II27705);
  nand NAND2_5439(WX9015,II27706,II27707);
  nand NAND2_5440(II27712,WX8395,CRC_OUT_3_5);
  nand NAND2_5441(II27713,WX8395,II27712);
  nand NAND2_5442(II27714,CRC_OUT_3_5,II27712);
  nand NAND2_5443(WX9016,II27713,II27714);
  nand NAND2_5444(II27719,WX8396,CRC_OUT_3_4);
  nand NAND2_5445(II27720,WX8396,II27719);
  nand NAND2_5446(II27721,CRC_OUT_3_4,II27719);
  nand NAND2_5447(WX9017,II27720,II27721);
  nand NAND2_5448(II27726,WX8398,CRC_OUT_3_2);
  nand NAND2_5449(II27727,WX8398,II27726);
  nand NAND2_5450(II27728,CRC_OUT_3_2,II27726);
  nand NAND2_5451(WX9018,II27727,II27728);
  nand NAND2_5452(II27733,WX8399,CRC_OUT_3_1);
  nand NAND2_5453(II27734,WX8399,II27733);
  nand NAND2_5454(II27735,CRC_OUT_3_1,II27733);
  nand NAND2_5455(WX9019,II27734,II27735);
  nand NAND2_5456(II27740,WX8400,CRC_OUT_3_0);
  nand NAND2_5457(II27741,WX8400,II27740);
  nand NAND2_5458(II27742,CRC_OUT_3_0,II27740);
  nand NAND2_5459(WX9020,II27741,II27742);
  nand NAND2_5460(II30023,WX10052,WX9696);
  nand NAND2_5461(II30024,WX10052,II30023);
  nand NAND2_5462(II30025,WX9696,II30023);
  nand NAND2_5463(II30022,II30024,II30025);
  nand NAND2_5464(II30030,WX9760,II30022);
  nand NAND2_5465(II30031,WX9760,II30030);
  nand NAND2_5466(II30032,II30022,II30030);
  nand NAND2_5467(II30021,II30031,II30032);
  nand NAND2_5468(II30038,WX9824,WX9888);
  nand NAND2_5469(II30039,WX9824,II30038);
  nand NAND2_5470(II30040,WX9888,II30038);
  nand NAND2_5471(II30037,II30039,II30040);
  nand NAND2_5472(II30045,II30021,II30037);
  nand NAND2_5473(II30046,II30021,II30045);
  nand NAND2_5474(II30047,II30037,II30045);
  nand NAND2_5475(WX9951,II30046,II30047);
  nand NAND2_5476(II30054,WX10052,WX9698);
  nand NAND2_5477(II30055,WX10052,II30054);
  nand NAND2_5478(II30056,WX9698,II30054);
  nand NAND2_5479(II30053,II30055,II30056);
  nand NAND2_5480(II30061,WX9762,II30053);
  nand NAND2_5481(II30062,WX9762,II30061);
  nand NAND2_5482(II30063,II30053,II30061);
  nand NAND2_5483(II30052,II30062,II30063);
  nand NAND2_5484(II30069,WX9826,WX9890);
  nand NAND2_5485(II30070,WX9826,II30069);
  nand NAND2_5486(II30071,WX9890,II30069);
  nand NAND2_5487(II30068,II30070,II30071);
  nand NAND2_5488(II30076,II30052,II30068);
  nand NAND2_5489(II30077,II30052,II30076);
  nand NAND2_5490(II30078,II30068,II30076);
  nand NAND2_5491(WX9952,II30077,II30078);
  nand NAND2_5492(II30085,WX10052,WX9700);
  nand NAND2_5493(II30086,WX10052,II30085);
  nand NAND2_5494(II30087,WX9700,II30085);
  nand NAND2_5495(II30084,II30086,II30087);
  nand NAND2_5496(II30092,WX9764,II30084);
  nand NAND2_5497(II30093,WX9764,II30092);
  nand NAND2_5498(II30094,II30084,II30092);
  nand NAND2_5499(II30083,II30093,II30094);
  nand NAND2_5500(II30100,WX9828,WX9892);
  nand NAND2_5501(II30101,WX9828,II30100);
  nand NAND2_5502(II30102,WX9892,II30100);
  nand NAND2_5503(II30099,II30101,II30102);
  nand NAND2_5504(II30107,II30083,II30099);
  nand NAND2_5505(II30108,II30083,II30107);
  nand NAND2_5506(II30109,II30099,II30107);
  nand NAND2_5507(WX9953,II30108,II30109);
  nand NAND2_5508(II30116,WX10052,WX9702);
  nand NAND2_5509(II30117,WX10052,II30116);
  nand NAND2_5510(II30118,WX9702,II30116);
  nand NAND2_5511(II30115,II30117,II30118);
  nand NAND2_5512(II30123,WX9766,II30115);
  nand NAND2_5513(II30124,WX9766,II30123);
  nand NAND2_5514(II30125,II30115,II30123);
  nand NAND2_5515(II30114,II30124,II30125);
  nand NAND2_5516(II30131,WX9830,WX9894);
  nand NAND2_5517(II30132,WX9830,II30131);
  nand NAND2_5518(II30133,WX9894,II30131);
  nand NAND2_5519(II30130,II30132,II30133);
  nand NAND2_5520(II30138,II30114,II30130);
  nand NAND2_5521(II30139,II30114,II30138);
  nand NAND2_5522(II30140,II30130,II30138);
  nand NAND2_5523(WX9954,II30139,II30140);
  nand NAND2_5524(II30147,WX10052,WX9704);
  nand NAND2_5525(II30148,WX10052,II30147);
  nand NAND2_5526(II30149,WX9704,II30147);
  nand NAND2_5527(II30146,II30148,II30149);
  nand NAND2_5528(II30154,WX9768,II30146);
  nand NAND2_5529(II30155,WX9768,II30154);
  nand NAND2_5530(II30156,II30146,II30154);
  nand NAND2_5531(II30145,II30155,II30156);
  nand NAND2_5532(II30162,WX9832,WX9896);
  nand NAND2_5533(II30163,WX9832,II30162);
  nand NAND2_5534(II30164,WX9896,II30162);
  nand NAND2_5535(II30161,II30163,II30164);
  nand NAND2_5536(II30169,II30145,II30161);
  nand NAND2_5537(II30170,II30145,II30169);
  nand NAND2_5538(II30171,II30161,II30169);
  nand NAND2_5539(WX9955,II30170,II30171);
  nand NAND2_5540(II30178,WX10052,WX9706);
  nand NAND2_5541(II30179,WX10052,II30178);
  nand NAND2_5542(II30180,WX9706,II30178);
  nand NAND2_5543(II30177,II30179,II30180);
  nand NAND2_5544(II30185,WX9770,II30177);
  nand NAND2_5545(II30186,WX9770,II30185);
  nand NAND2_5546(II30187,II30177,II30185);
  nand NAND2_5547(II30176,II30186,II30187);
  nand NAND2_5548(II30193,WX9834,WX9898);
  nand NAND2_5549(II30194,WX9834,II30193);
  nand NAND2_5550(II30195,WX9898,II30193);
  nand NAND2_5551(II30192,II30194,II30195);
  nand NAND2_5552(II30200,II30176,II30192);
  nand NAND2_5553(II30201,II30176,II30200);
  nand NAND2_5554(II30202,II30192,II30200);
  nand NAND2_5555(WX9956,II30201,II30202);
  nand NAND2_5556(II30209,WX10052,WX9708);
  nand NAND2_5557(II30210,WX10052,II30209);
  nand NAND2_5558(II30211,WX9708,II30209);
  nand NAND2_5559(II30208,II30210,II30211);
  nand NAND2_5560(II30216,WX9772,II30208);
  nand NAND2_5561(II30217,WX9772,II30216);
  nand NAND2_5562(II30218,II30208,II30216);
  nand NAND2_5563(II30207,II30217,II30218);
  nand NAND2_5564(II30224,WX9836,WX9900);
  nand NAND2_5565(II30225,WX9836,II30224);
  nand NAND2_5566(II30226,WX9900,II30224);
  nand NAND2_5567(II30223,II30225,II30226);
  nand NAND2_5568(II30231,II30207,II30223);
  nand NAND2_5569(II30232,II30207,II30231);
  nand NAND2_5570(II30233,II30223,II30231);
  nand NAND2_5571(WX9957,II30232,II30233);
  nand NAND2_5572(II30240,WX10052,WX9710);
  nand NAND2_5573(II30241,WX10052,II30240);
  nand NAND2_5574(II30242,WX9710,II30240);
  nand NAND2_5575(II30239,II30241,II30242);
  nand NAND2_5576(II30247,WX9774,II30239);
  nand NAND2_5577(II30248,WX9774,II30247);
  nand NAND2_5578(II30249,II30239,II30247);
  nand NAND2_5579(II30238,II30248,II30249);
  nand NAND2_5580(II30255,WX9838,WX9902);
  nand NAND2_5581(II30256,WX9838,II30255);
  nand NAND2_5582(II30257,WX9902,II30255);
  nand NAND2_5583(II30254,II30256,II30257);
  nand NAND2_5584(II30262,II30238,II30254);
  nand NAND2_5585(II30263,II30238,II30262);
  nand NAND2_5586(II30264,II30254,II30262);
  nand NAND2_5587(WX9958,II30263,II30264);
  nand NAND2_5588(II30271,WX10052,WX9712);
  nand NAND2_5589(II30272,WX10052,II30271);
  nand NAND2_5590(II30273,WX9712,II30271);
  nand NAND2_5591(II30270,II30272,II30273);
  nand NAND2_5592(II30278,WX9776,II30270);
  nand NAND2_5593(II30279,WX9776,II30278);
  nand NAND2_5594(II30280,II30270,II30278);
  nand NAND2_5595(II30269,II30279,II30280);
  nand NAND2_5596(II30286,WX9840,WX9904);
  nand NAND2_5597(II30287,WX9840,II30286);
  nand NAND2_5598(II30288,WX9904,II30286);
  nand NAND2_5599(II30285,II30287,II30288);
  nand NAND2_5600(II30293,II30269,II30285);
  nand NAND2_5601(II30294,II30269,II30293);
  nand NAND2_5602(II30295,II30285,II30293);
  nand NAND2_5603(WX9959,II30294,II30295);
  nand NAND2_5604(II30302,WX10052,WX9714);
  nand NAND2_5605(II30303,WX10052,II30302);
  nand NAND2_5606(II30304,WX9714,II30302);
  nand NAND2_5607(II30301,II30303,II30304);
  nand NAND2_5608(II30309,WX9778,II30301);
  nand NAND2_5609(II30310,WX9778,II30309);
  nand NAND2_5610(II30311,II30301,II30309);
  nand NAND2_5611(II30300,II30310,II30311);
  nand NAND2_5612(II30317,WX9842,WX9906);
  nand NAND2_5613(II30318,WX9842,II30317);
  nand NAND2_5614(II30319,WX9906,II30317);
  nand NAND2_5615(II30316,II30318,II30319);
  nand NAND2_5616(II30324,II30300,II30316);
  nand NAND2_5617(II30325,II30300,II30324);
  nand NAND2_5618(II30326,II30316,II30324);
  nand NAND2_5619(WX9960,II30325,II30326);
  nand NAND2_5620(II30333,WX10052,WX9716);
  nand NAND2_5621(II30334,WX10052,II30333);
  nand NAND2_5622(II30335,WX9716,II30333);
  nand NAND2_5623(II30332,II30334,II30335);
  nand NAND2_5624(II30340,WX9780,II30332);
  nand NAND2_5625(II30341,WX9780,II30340);
  nand NAND2_5626(II30342,II30332,II30340);
  nand NAND2_5627(II30331,II30341,II30342);
  nand NAND2_5628(II30348,WX9844,WX9908);
  nand NAND2_5629(II30349,WX9844,II30348);
  nand NAND2_5630(II30350,WX9908,II30348);
  nand NAND2_5631(II30347,II30349,II30350);
  nand NAND2_5632(II30355,II30331,II30347);
  nand NAND2_5633(II30356,II30331,II30355);
  nand NAND2_5634(II30357,II30347,II30355);
  nand NAND2_5635(WX9961,II30356,II30357);
  nand NAND2_5636(II30364,WX10052,WX9718);
  nand NAND2_5637(II30365,WX10052,II30364);
  nand NAND2_5638(II30366,WX9718,II30364);
  nand NAND2_5639(II30363,II30365,II30366);
  nand NAND2_5640(II30371,WX9782,II30363);
  nand NAND2_5641(II30372,WX9782,II30371);
  nand NAND2_5642(II30373,II30363,II30371);
  nand NAND2_5643(II30362,II30372,II30373);
  nand NAND2_5644(II30379,WX9846,WX9910);
  nand NAND2_5645(II30380,WX9846,II30379);
  nand NAND2_5646(II30381,WX9910,II30379);
  nand NAND2_5647(II30378,II30380,II30381);
  nand NAND2_5648(II30386,II30362,II30378);
  nand NAND2_5649(II30387,II30362,II30386);
  nand NAND2_5650(II30388,II30378,II30386);
  nand NAND2_5651(WX9962,II30387,II30388);
  nand NAND2_5652(II30395,WX10052,WX9720);
  nand NAND2_5653(II30396,WX10052,II30395);
  nand NAND2_5654(II30397,WX9720,II30395);
  nand NAND2_5655(II30394,II30396,II30397);
  nand NAND2_5656(II30402,WX9784,II30394);
  nand NAND2_5657(II30403,WX9784,II30402);
  nand NAND2_5658(II30404,II30394,II30402);
  nand NAND2_5659(II30393,II30403,II30404);
  nand NAND2_5660(II30410,WX9848,WX9912);
  nand NAND2_5661(II30411,WX9848,II30410);
  nand NAND2_5662(II30412,WX9912,II30410);
  nand NAND2_5663(II30409,II30411,II30412);
  nand NAND2_5664(II30417,II30393,II30409);
  nand NAND2_5665(II30418,II30393,II30417);
  nand NAND2_5666(II30419,II30409,II30417);
  nand NAND2_5667(WX9963,II30418,II30419);
  nand NAND2_5668(II30426,WX10052,WX9722);
  nand NAND2_5669(II30427,WX10052,II30426);
  nand NAND2_5670(II30428,WX9722,II30426);
  nand NAND2_5671(II30425,II30427,II30428);
  nand NAND2_5672(II30433,WX9786,II30425);
  nand NAND2_5673(II30434,WX9786,II30433);
  nand NAND2_5674(II30435,II30425,II30433);
  nand NAND2_5675(II30424,II30434,II30435);
  nand NAND2_5676(II30441,WX9850,WX9914);
  nand NAND2_5677(II30442,WX9850,II30441);
  nand NAND2_5678(II30443,WX9914,II30441);
  nand NAND2_5679(II30440,II30442,II30443);
  nand NAND2_5680(II30448,II30424,II30440);
  nand NAND2_5681(II30449,II30424,II30448);
  nand NAND2_5682(II30450,II30440,II30448);
  nand NAND2_5683(WX9964,II30449,II30450);
  nand NAND2_5684(II30457,WX10052,WX9724);
  nand NAND2_5685(II30458,WX10052,II30457);
  nand NAND2_5686(II30459,WX9724,II30457);
  nand NAND2_5687(II30456,II30458,II30459);
  nand NAND2_5688(II30464,WX9788,II30456);
  nand NAND2_5689(II30465,WX9788,II30464);
  nand NAND2_5690(II30466,II30456,II30464);
  nand NAND2_5691(II30455,II30465,II30466);
  nand NAND2_5692(II30472,WX9852,WX9916);
  nand NAND2_5693(II30473,WX9852,II30472);
  nand NAND2_5694(II30474,WX9916,II30472);
  nand NAND2_5695(II30471,II30473,II30474);
  nand NAND2_5696(II30479,II30455,II30471);
  nand NAND2_5697(II30480,II30455,II30479);
  nand NAND2_5698(II30481,II30471,II30479);
  nand NAND2_5699(WX9965,II30480,II30481);
  nand NAND2_5700(II30488,WX10052,WX9726);
  nand NAND2_5701(II30489,WX10052,II30488);
  nand NAND2_5702(II30490,WX9726,II30488);
  nand NAND2_5703(II30487,II30489,II30490);
  nand NAND2_5704(II30495,WX9790,II30487);
  nand NAND2_5705(II30496,WX9790,II30495);
  nand NAND2_5706(II30497,II30487,II30495);
  nand NAND2_5707(II30486,II30496,II30497);
  nand NAND2_5708(II30503,WX9854,WX9918);
  nand NAND2_5709(II30504,WX9854,II30503);
  nand NAND2_5710(II30505,WX9918,II30503);
  nand NAND2_5711(II30502,II30504,II30505);
  nand NAND2_5712(II30510,II30486,II30502);
  nand NAND2_5713(II30511,II30486,II30510);
  nand NAND2_5714(II30512,II30502,II30510);
  nand NAND2_5715(WX9966,II30511,II30512);
  nand NAND2_5716(II30519,WX10053,WX9728);
  nand NAND2_5717(II30520,WX10053,II30519);
  nand NAND2_5718(II30521,WX9728,II30519);
  nand NAND2_5719(II30518,II30520,II30521);
  nand NAND2_5720(II30526,WX9792,II30518);
  nand NAND2_5721(II30527,WX9792,II30526);
  nand NAND2_5722(II30528,II30518,II30526);
  nand NAND2_5723(II30517,II30527,II30528);
  nand NAND2_5724(II30534,WX9856,WX9920);
  nand NAND2_5725(II30535,WX9856,II30534);
  nand NAND2_5726(II30536,WX9920,II30534);
  nand NAND2_5727(II30533,II30535,II30536);
  nand NAND2_5728(II30541,II30517,II30533);
  nand NAND2_5729(II30542,II30517,II30541);
  nand NAND2_5730(II30543,II30533,II30541);
  nand NAND2_5731(WX9967,II30542,II30543);
  nand NAND2_5732(II30550,WX10053,WX9730);
  nand NAND2_5733(II30551,WX10053,II30550);
  nand NAND2_5734(II30552,WX9730,II30550);
  nand NAND2_5735(II30549,II30551,II30552);
  nand NAND2_5736(II30557,WX9794,II30549);
  nand NAND2_5737(II30558,WX9794,II30557);
  nand NAND2_5738(II30559,II30549,II30557);
  nand NAND2_5739(II30548,II30558,II30559);
  nand NAND2_5740(II30565,WX9858,WX9922);
  nand NAND2_5741(II30566,WX9858,II30565);
  nand NAND2_5742(II30567,WX9922,II30565);
  nand NAND2_5743(II30564,II30566,II30567);
  nand NAND2_5744(II30572,II30548,II30564);
  nand NAND2_5745(II30573,II30548,II30572);
  nand NAND2_5746(II30574,II30564,II30572);
  nand NAND2_5747(WX9968,II30573,II30574);
  nand NAND2_5748(II30581,WX10053,WX9732);
  nand NAND2_5749(II30582,WX10053,II30581);
  nand NAND2_5750(II30583,WX9732,II30581);
  nand NAND2_5751(II30580,II30582,II30583);
  nand NAND2_5752(II30588,WX9796,II30580);
  nand NAND2_5753(II30589,WX9796,II30588);
  nand NAND2_5754(II30590,II30580,II30588);
  nand NAND2_5755(II30579,II30589,II30590);
  nand NAND2_5756(II30596,WX9860,WX9924);
  nand NAND2_5757(II30597,WX9860,II30596);
  nand NAND2_5758(II30598,WX9924,II30596);
  nand NAND2_5759(II30595,II30597,II30598);
  nand NAND2_5760(II30603,II30579,II30595);
  nand NAND2_5761(II30604,II30579,II30603);
  nand NAND2_5762(II30605,II30595,II30603);
  nand NAND2_5763(WX9969,II30604,II30605);
  nand NAND2_5764(II30612,WX10053,WX9734);
  nand NAND2_5765(II30613,WX10053,II30612);
  nand NAND2_5766(II30614,WX9734,II30612);
  nand NAND2_5767(II30611,II30613,II30614);
  nand NAND2_5768(II30619,WX9798,II30611);
  nand NAND2_5769(II30620,WX9798,II30619);
  nand NAND2_5770(II30621,II30611,II30619);
  nand NAND2_5771(II30610,II30620,II30621);
  nand NAND2_5772(II30627,WX9862,WX9926);
  nand NAND2_5773(II30628,WX9862,II30627);
  nand NAND2_5774(II30629,WX9926,II30627);
  nand NAND2_5775(II30626,II30628,II30629);
  nand NAND2_5776(II30634,II30610,II30626);
  nand NAND2_5777(II30635,II30610,II30634);
  nand NAND2_5778(II30636,II30626,II30634);
  nand NAND2_5779(WX9970,II30635,II30636);
  nand NAND2_5780(II30643,WX10053,WX9736);
  nand NAND2_5781(II30644,WX10053,II30643);
  nand NAND2_5782(II30645,WX9736,II30643);
  nand NAND2_5783(II30642,II30644,II30645);
  nand NAND2_5784(II30650,WX9800,II30642);
  nand NAND2_5785(II30651,WX9800,II30650);
  nand NAND2_5786(II30652,II30642,II30650);
  nand NAND2_5787(II30641,II30651,II30652);
  nand NAND2_5788(II30658,WX9864,WX9928);
  nand NAND2_5789(II30659,WX9864,II30658);
  nand NAND2_5790(II30660,WX9928,II30658);
  nand NAND2_5791(II30657,II30659,II30660);
  nand NAND2_5792(II30665,II30641,II30657);
  nand NAND2_5793(II30666,II30641,II30665);
  nand NAND2_5794(II30667,II30657,II30665);
  nand NAND2_5795(WX9971,II30666,II30667);
  nand NAND2_5796(II30674,WX10053,WX9738);
  nand NAND2_5797(II30675,WX10053,II30674);
  nand NAND2_5798(II30676,WX9738,II30674);
  nand NAND2_5799(II30673,II30675,II30676);
  nand NAND2_5800(II30681,WX9802,II30673);
  nand NAND2_5801(II30682,WX9802,II30681);
  nand NAND2_5802(II30683,II30673,II30681);
  nand NAND2_5803(II30672,II30682,II30683);
  nand NAND2_5804(II30689,WX9866,WX9930);
  nand NAND2_5805(II30690,WX9866,II30689);
  nand NAND2_5806(II30691,WX9930,II30689);
  nand NAND2_5807(II30688,II30690,II30691);
  nand NAND2_5808(II30696,II30672,II30688);
  nand NAND2_5809(II30697,II30672,II30696);
  nand NAND2_5810(II30698,II30688,II30696);
  nand NAND2_5811(WX9972,II30697,II30698);
  nand NAND2_5812(II30705,WX10053,WX9740);
  nand NAND2_5813(II30706,WX10053,II30705);
  nand NAND2_5814(II30707,WX9740,II30705);
  nand NAND2_5815(II30704,II30706,II30707);
  nand NAND2_5816(II30712,WX9804,II30704);
  nand NAND2_5817(II30713,WX9804,II30712);
  nand NAND2_5818(II30714,II30704,II30712);
  nand NAND2_5819(II30703,II30713,II30714);
  nand NAND2_5820(II30720,WX9868,WX9932);
  nand NAND2_5821(II30721,WX9868,II30720);
  nand NAND2_5822(II30722,WX9932,II30720);
  nand NAND2_5823(II30719,II30721,II30722);
  nand NAND2_5824(II30727,II30703,II30719);
  nand NAND2_5825(II30728,II30703,II30727);
  nand NAND2_5826(II30729,II30719,II30727);
  nand NAND2_5827(WX9973,II30728,II30729);
  nand NAND2_5828(II30736,WX10053,WX9742);
  nand NAND2_5829(II30737,WX10053,II30736);
  nand NAND2_5830(II30738,WX9742,II30736);
  nand NAND2_5831(II30735,II30737,II30738);
  nand NAND2_5832(II30743,WX9806,II30735);
  nand NAND2_5833(II30744,WX9806,II30743);
  nand NAND2_5834(II30745,II30735,II30743);
  nand NAND2_5835(II30734,II30744,II30745);
  nand NAND2_5836(II30751,WX9870,WX9934);
  nand NAND2_5837(II30752,WX9870,II30751);
  nand NAND2_5838(II30753,WX9934,II30751);
  nand NAND2_5839(II30750,II30752,II30753);
  nand NAND2_5840(II30758,II30734,II30750);
  nand NAND2_5841(II30759,II30734,II30758);
  nand NAND2_5842(II30760,II30750,II30758);
  nand NAND2_5843(WX9974,II30759,II30760);
  nand NAND2_5844(II30767,WX10053,WX9744);
  nand NAND2_5845(II30768,WX10053,II30767);
  nand NAND2_5846(II30769,WX9744,II30767);
  nand NAND2_5847(II30766,II30768,II30769);
  nand NAND2_5848(II30774,WX9808,II30766);
  nand NAND2_5849(II30775,WX9808,II30774);
  nand NAND2_5850(II30776,II30766,II30774);
  nand NAND2_5851(II30765,II30775,II30776);
  nand NAND2_5852(II30782,WX9872,WX9936);
  nand NAND2_5853(II30783,WX9872,II30782);
  nand NAND2_5854(II30784,WX9936,II30782);
  nand NAND2_5855(II30781,II30783,II30784);
  nand NAND2_5856(II30789,II30765,II30781);
  nand NAND2_5857(II30790,II30765,II30789);
  nand NAND2_5858(II30791,II30781,II30789);
  nand NAND2_5859(WX9975,II30790,II30791);
  nand NAND2_5860(II30798,WX10053,WX9746);
  nand NAND2_5861(II30799,WX10053,II30798);
  nand NAND2_5862(II30800,WX9746,II30798);
  nand NAND2_5863(II30797,II30799,II30800);
  nand NAND2_5864(II30805,WX9810,II30797);
  nand NAND2_5865(II30806,WX9810,II30805);
  nand NAND2_5866(II30807,II30797,II30805);
  nand NAND2_5867(II30796,II30806,II30807);
  nand NAND2_5868(II30813,WX9874,WX9938);
  nand NAND2_5869(II30814,WX9874,II30813);
  nand NAND2_5870(II30815,WX9938,II30813);
  nand NAND2_5871(II30812,II30814,II30815);
  nand NAND2_5872(II30820,II30796,II30812);
  nand NAND2_5873(II30821,II30796,II30820);
  nand NAND2_5874(II30822,II30812,II30820);
  nand NAND2_5875(WX9976,II30821,II30822);
  nand NAND2_5876(II30829,WX10053,WX9748);
  nand NAND2_5877(II30830,WX10053,II30829);
  nand NAND2_5878(II30831,WX9748,II30829);
  nand NAND2_5879(II30828,II30830,II30831);
  nand NAND2_5880(II30836,WX9812,II30828);
  nand NAND2_5881(II30837,WX9812,II30836);
  nand NAND2_5882(II30838,II30828,II30836);
  nand NAND2_5883(II30827,II30837,II30838);
  nand NAND2_5884(II30844,WX9876,WX9940);
  nand NAND2_5885(II30845,WX9876,II30844);
  nand NAND2_5886(II30846,WX9940,II30844);
  nand NAND2_5887(II30843,II30845,II30846);
  nand NAND2_5888(II30851,II30827,II30843);
  nand NAND2_5889(II30852,II30827,II30851);
  nand NAND2_5890(II30853,II30843,II30851);
  nand NAND2_5891(WX9977,II30852,II30853);
  nand NAND2_5892(II30860,WX10053,WX9750);
  nand NAND2_5893(II30861,WX10053,II30860);
  nand NAND2_5894(II30862,WX9750,II30860);
  nand NAND2_5895(II30859,II30861,II30862);
  nand NAND2_5896(II30867,WX9814,II30859);
  nand NAND2_5897(II30868,WX9814,II30867);
  nand NAND2_5898(II30869,II30859,II30867);
  nand NAND2_5899(II30858,II30868,II30869);
  nand NAND2_5900(II30875,WX9878,WX9942);
  nand NAND2_5901(II30876,WX9878,II30875);
  nand NAND2_5902(II30877,WX9942,II30875);
  nand NAND2_5903(II30874,II30876,II30877);
  nand NAND2_5904(II30882,II30858,II30874);
  nand NAND2_5905(II30883,II30858,II30882);
  nand NAND2_5906(II30884,II30874,II30882);
  nand NAND2_5907(WX9978,II30883,II30884);
  nand NAND2_5908(II30891,WX10053,WX9752);
  nand NAND2_5909(II30892,WX10053,II30891);
  nand NAND2_5910(II30893,WX9752,II30891);
  nand NAND2_5911(II30890,II30892,II30893);
  nand NAND2_5912(II30898,WX9816,II30890);
  nand NAND2_5913(II30899,WX9816,II30898);
  nand NAND2_5914(II30900,II30890,II30898);
  nand NAND2_5915(II30889,II30899,II30900);
  nand NAND2_5916(II30906,WX9880,WX9944);
  nand NAND2_5917(II30907,WX9880,II30906);
  nand NAND2_5918(II30908,WX9944,II30906);
  nand NAND2_5919(II30905,II30907,II30908);
  nand NAND2_5920(II30913,II30889,II30905);
  nand NAND2_5921(II30914,II30889,II30913);
  nand NAND2_5922(II30915,II30905,II30913);
  nand NAND2_5923(WX9979,II30914,II30915);
  nand NAND2_5924(II30922,WX10053,WX9754);
  nand NAND2_5925(II30923,WX10053,II30922);
  nand NAND2_5926(II30924,WX9754,II30922);
  nand NAND2_5927(II30921,II30923,II30924);
  nand NAND2_5928(II30929,WX9818,II30921);
  nand NAND2_5929(II30930,WX9818,II30929);
  nand NAND2_5930(II30931,II30921,II30929);
  nand NAND2_5931(II30920,II30930,II30931);
  nand NAND2_5932(II30937,WX9882,WX9946);
  nand NAND2_5933(II30938,WX9882,II30937);
  nand NAND2_5934(II30939,WX9946,II30937);
  nand NAND2_5935(II30936,II30938,II30939);
  nand NAND2_5936(II30944,II30920,II30936);
  nand NAND2_5937(II30945,II30920,II30944);
  nand NAND2_5938(II30946,II30936,II30944);
  nand NAND2_5939(WX9980,II30945,II30946);
  nand NAND2_5940(II30953,WX10053,WX9756);
  nand NAND2_5941(II30954,WX10053,II30953);
  nand NAND2_5942(II30955,WX9756,II30953);
  nand NAND2_5943(II30952,II30954,II30955);
  nand NAND2_5944(II30960,WX9820,II30952);
  nand NAND2_5945(II30961,WX9820,II30960);
  nand NAND2_5946(II30962,II30952,II30960);
  nand NAND2_5947(II30951,II30961,II30962);
  nand NAND2_5948(II30968,WX9884,WX9948);
  nand NAND2_5949(II30969,WX9884,II30968);
  nand NAND2_5950(II30970,WX9948,II30968);
  nand NAND2_5951(II30967,II30969,II30970);
  nand NAND2_5952(II30975,II30951,II30967);
  nand NAND2_5953(II30976,II30951,II30975);
  nand NAND2_5954(II30977,II30967,II30975);
  nand NAND2_5955(WX9981,II30976,II30977);
  nand NAND2_5956(II30984,WX10053,WX9758);
  nand NAND2_5957(II30985,WX10053,II30984);
  nand NAND2_5958(II30986,WX9758,II30984);
  nand NAND2_5959(II30983,II30985,II30986);
  nand NAND2_5960(II30991,WX9822,II30983);
  nand NAND2_5961(II30992,WX9822,II30991);
  nand NAND2_5962(II30993,II30983,II30991);
  nand NAND2_5963(II30982,II30992,II30993);
  nand NAND2_5964(II30999,WX9886,WX9950);
  nand NAND2_5965(II31000,WX9886,II30999);
  nand NAND2_5966(II31001,WX9950,II30999);
  nand NAND2_5967(II30998,II31000,II31001);
  nand NAND2_5968(II31006,II30982,II30998);
  nand NAND2_5969(II31007,II30982,II31006);
  nand NAND2_5970(II31008,II30998,II31006);
  nand NAND2_5971(WX9982,II31007,II31008);
  nand NAND2_5972(II31087,WX9631,WX9536);
  nand NAND2_5973(II31088,WX9631,II31087);
  nand NAND2_5974(II31089,WX9536,II31087);
  nand NAND2_5975(WX10057,II31088,II31089);
  nand NAND2_5976(II31100,WX9632,WX9538);
  nand NAND2_5977(II31101,WX9632,II31100);
  nand NAND2_5978(II31102,WX9538,II31100);
  nand NAND2_5979(WX10064,II31101,II31102);
  nand NAND2_5980(II31113,WX9633,WX9540);
  nand NAND2_5981(II31114,WX9633,II31113);
  nand NAND2_5982(II31115,WX9540,II31113);
  nand NAND2_5983(WX10071,II31114,II31115);
  nand NAND2_5984(II31126,WX9634,WX9542);
  nand NAND2_5985(II31127,WX9634,II31126);
  nand NAND2_5986(II31128,WX9542,II31126);
  nand NAND2_5987(WX10078,II31127,II31128);
  nand NAND2_5988(II31139,WX9635,WX9544);
  nand NAND2_5989(II31140,WX9635,II31139);
  nand NAND2_5990(II31141,WX9544,II31139);
  nand NAND2_5991(WX10085,II31140,II31141);
  nand NAND2_5992(II31152,WX9636,WX9546);
  nand NAND2_5993(II31153,WX9636,II31152);
  nand NAND2_5994(II31154,WX9546,II31152);
  nand NAND2_5995(WX10092,II31153,II31154);
  nand NAND2_5996(II31165,WX9637,WX9548);
  nand NAND2_5997(II31166,WX9637,II31165);
  nand NAND2_5998(II31167,WX9548,II31165);
  nand NAND2_5999(WX10099,II31166,II31167);
  nand NAND2_6000(II31178,WX9638,WX9550);
  nand NAND2_6001(II31179,WX9638,II31178);
  nand NAND2_6002(II31180,WX9550,II31178);
  nand NAND2_6003(WX10106,II31179,II31180);
  nand NAND2_6004(II31191,WX9639,WX9552);
  nand NAND2_6005(II31192,WX9639,II31191);
  nand NAND2_6006(II31193,WX9552,II31191);
  nand NAND2_6007(WX10113,II31192,II31193);
  nand NAND2_6008(II31204,WX9640,WX9554);
  nand NAND2_6009(II31205,WX9640,II31204);
  nand NAND2_6010(II31206,WX9554,II31204);
  nand NAND2_6011(WX10120,II31205,II31206);
  nand NAND2_6012(II31217,WX9641,WX9556);
  nand NAND2_6013(II31218,WX9641,II31217);
  nand NAND2_6014(II31219,WX9556,II31217);
  nand NAND2_6015(WX10127,II31218,II31219);
  nand NAND2_6016(II31230,WX9642,WX9558);
  nand NAND2_6017(II31231,WX9642,II31230);
  nand NAND2_6018(II31232,WX9558,II31230);
  nand NAND2_6019(WX10134,II31231,II31232);
  nand NAND2_6020(II31243,WX9643,WX9560);
  nand NAND2_6021(II31244,WX9643,II31243);
  nand NAND2_6022(II31245,WX9560,II31243);
  nand NAND2_6023(WX10141,II31244,II31245);
  nand NAND2_6024(II31256,WX9644,WX9562);
  nand NAND2_6025(II31257,WX9644,II31256);
  nand NAND2_6026(II31258,WX9562,II31256);
  nand NAND2_6027(WX10148,II31257,II31258);
  nand NAND2_6028(II31269,WX9645,WX9564);
  nand NAND2_6029(II31270,WX9645,II31269);
  nand NAND2_6030(II31271,WX9564,II31269);
  nand NAND2_6031(WX10155,II31270,II31271);
  nand NAND2_6032(II31282,WX9646,WX9566);
  nand NAND2_6033(II31283,WX9646,II31282);
  nand NAND2_6034(II31284,WX9566,II31282);
  nand NAND2_6035(WX10162,II31283,II31284);
  nand NAND2_6036(II31295,WX9647,WX9568);
  nand NAND2_6037(II31296,WX9647,II31295);
  nand NAND2_6038(II31297,WX9568,II31295);
  nand NAND2_6039(WX10169,II31296,II31297);
  nand NAND2_6040(II31308,WX9648,WX9570);
  nand NAND2_6041(II31309,WX9648,II31308);
  nand NAND2_6042(II31310,WX9570,II31308);
  nand NAND2_6043(WX10176,II31309,II31310);
  nand NAND2_6044(II31321,WX9649,WX9572);
  nand NAND2_6045(II31322,WX9649,II31321);
  nand NAND2_6046(II31323,WX9572,II31321);
  nand NAND2_6047(WX10183,II31322,II31323);
  nand NAND2_6048(II31334,WX9650,WX9574);
  nand NAND2_6049(II31335,WX9650,II31334);
  nand NAND2_6050(II31336,WX9574,II31334);
  nand NAND2_6051(WX10190,II31335,II31336);
  nand NAND2_6052(II31347,WX9651,WX9576);
  nand NAND2_6053(II31348,WX9651,II31347);
  nand NAND2_6054(II31349,WX9576,II31347);
  nand NAND2_6055(WX10197,II31348,II31349);
  nand NAND2_6056(II31360,WX9652,WX9578);
  nand NAND2_6057(II31361,WX9652,II31360);
  nand NAND2_6058(II31362,WX9578,II31360);
  nand NAND2_6059(WX10204,II31361,II31362);
  nand NAND2_6060(II31373,WX9653,WX9580);
  nand NAND2_6061(II31374,WX9653,II31373);
  nand NAND2_6062(II31375,WX9580,II31373);
  nand NAND2_6063(WX10211,II31374,II31375);
  nand NAND2_6064(II31386,WX9654,WX9582);
  nand NAND2_6065(II31387,WX9654,II31386);
  nand NAND2_6066(II31388,WX9582,II31386);
  nand NAND2_6067(WX10218,II31387,II31388);
  nand NAND2_6068(II31399,WX9655,WX9584);
  nand NAND2_6069(II31400,WX9655,II31399);
  nand NAND2_6070(II31401,WX9584,II31399);
  nand NAND2_6071(WX10225,II31400,II31401);
  nand NAND2_6072(II31412,WX9656,WX9586);
  nand NAND2_6073(II31413,WX9656,II31412);
  nand NAND2_6074(II31414,WX9586,II31412);
  nand NAND2_6075(WX10232,II31413,II31414);
  nand NAND2_6076(II31425,WX9657,WX9588);
  nand NAND2_6077(II31426,WX9657,II31425);
  nand NAND2_6078(II31427,WX9588,II31425);
  nand NAND2_6079(WX10239,II31426,II31427);
  nand NAND2_6080(II31438,WX9658,WX9590);
  nand NAND2_6081(II31439,WX9658,II31438);
  nand NAND2_6082(II31440,WX9590,II31438);
  nand NAND2_6083(WX10246,II31439,II31440);
  nand NAND2_6084(II31451,WX9659,WX9592);
  nand NAND2_6085(II31452,WX9659,II31451);
  nand NAND2_6086(II31453,WX9592,II31451);
  nand NAND2_6087(WX10253,II31452,II31453);
  nand NAND2_6088(II31464,WX9660,WX9594);
  nand NAND2_6089(II31465,WX9660,II31464);
  nand NAND2_6090(II31466,WX9594,II31464);
  nand NAND2_6091(WX10260,II31465,II31466);
  nand NAND2_6092(II31477,WX9661,WX9596);
  nand NAND2_6093(II31478,WX9661,II31477);
  nand NAND2_6094(II31479,WX9596,II31477);
  nand NAND2_6095(WX10267,II31478,II31479);
  nand NAND2_6096(II31490,WX9662,WX9598);
  nand NAND2_6097(II31491,WX9662,II31490);
  nand NAND2_6098(II31492,WX9598,II31490);
  nand NAND2_6099(WX10274,II31491,II31492);
  nand NAND2_6100(II31505,WX9678,CRC_OUT_2_31);
  nand NAND2_6101(II31506,WX9678,II31505);
  nand NAND2_6102(II31507,CRC_OUT_2_31,II31505);
  nand NAND2_6103(II31504,II31506,II31507);
  nand NAND2_6104(II31512,CRC_OUT_2_15,II31504);
  nand NAND2_6105(II31513,CRC_OUT_2_15,II31512);
  nand NAND2_6106(II31514,II31504,II31512);
  nand NAND2_6107(WX10282,II31513,II31514);
  nand NAND2_6108(II31520,WX9683,CRC_OUT_2_31);
  nand NAND2_6109(II31521,WX9683,II31520);
  nand NAND2_6110(II31522,CRC_OUT_2_31,II31520);
  nand NAND2_6111(II31519,II31521,II31522);
  nand NAND2_6112(II31527,CRC_OUT_2_10,II31519);
  nand NAND2_6113(II31528,CRC_OUT_2_10,II31527);
  nand NAND2_6114(II31529,II31519,II31527);
  nand NAND2_6115(WX10283,II31528,II31529);
  nand NAND2_6116(II31535,WX9690,CRC_OUT_2_31);
  nand NAND2_6117(II31536,WX9690,II31535);
  nand NAND2_6118(II31537,CRC_OUT_2_31,II31535);
  nand NAND2_6119(II31534,II31536,II31537);
  nand NAND2_6120(II31542,CRC_OUT_2_3,II31534);
  nand NAND2_6121(II31543,CRC_OUT_2_3,II31542);
  nand NAND2_6122(II31544,II31534,II31542);
  nand NAND2_6123(WX10284,II31543,II31544);
  nand NAND2_6124(II31549,WX9694,CRC_OUT_2_31);
  nand NAND2_6125(II31550,WX9694,II31549);
  nand NAND2_6126(II31551,CRC_OUT_2_31,II31549);
  nand NAND2_6127(WX10285,II31550,II31551);
  nand NAND2_6128(II31556,WX9663,CRC_OUT_2_30);
  nand NAND2_6129(II31557,WX9663,II31556);
  nand NAND2_6130(II31558,CRC_OUT_2_30,II31556);
  nand NAND2_6131(WX10286,II31557,II31558);
  nand NAND2_6132(II31563,WX9664,CRC_OUT_2_29);
  nand NAND2_6133(II31564,WX9664,II31563);
  nand NAND2_6134(II31565,CRC_OUT_2_29,II31563);
  nand NAND2_6135(WX10287,II31564,II31565);
  nand NAND2_6136(II31570,WX9665,CRC_OUT_2_28);
  nand NAND2_6137(II31571,WX9665,II31570);
  nand NAND2_6138(II31572,CRC_OUT_2_28,II31570);
  nand NAND2_6139(WX10288,II31571,II31572);
  nand NAND2_6140(II31577,WX9666,CRC_OUT_2_27);
  nand NAND2_6141(II31578,WX9666,II31577);
  nand NAND2_6142(II31579,CRC_OUT_2_27,II31577);
  nand NAND2_6143(WX10289,II31578,II31579);
  nand NAND2_6144(II31584,WX9667,CRC_OUT_2_26);
  nand NAND2_6145(II31585,WX9667,II31584);
  nand NAND2_6146(II31586,CRC_OUT_2_26,II31584);
  nand NAND2_6147(WX10290,II31585,II31586);
  nand NAND2_6148(II31591,WX9668,CRC_OUT_2_25);
  nand NAND2_6149(II31592,WX9668,II31591);
  nand NAND2_6150(II31593,CRC_OUT_2_25,II31591);
  nand NAND2_6151(WX10291,II31592,II31593);
  nand NAND2_6152(II31598,WX9669,CRC_OUT_2_24);
  nand NAND2_6153(II31599,WX9669,II31598);
  nand NAND2_6154(II31600,CRC_OUT_2_24,II31598);
  nand NAND2_6155(WX10292,II31599,II31600);
  nand NAND2_6156(II31605,WX9670,CRC_OUT_2_23);
  nand NAND2_6157(II31606,WX9670,II31605);
  nand NAND2_6158(II31607,CRC_OUT_2_23,II31605);
  nand NAND2_6159(WX10293,II31606,II31607);
  nand NAND2_6160(II31612,WX9671,CRC_OUT_2_22);
  nand NAND2_6161(II31613,WX9671,II31612);
  nand NAND2_6162(II31614,CRC_OUT_2_22,II31612);
  nand NAND2_6163(WX10294,II31613,II31614);
  nand NAND2_6164(II31619,WX9672,CRC_OUT_2_21);
  nand NAND2_6165(II31620,WX9672,II31619);
  nand NAND2_6166(II31621,CRC_OUT_2_21,II31619);
  nand NAND2_6167(WX10295,II31620,II31621);
  nand NAND2_6168(II31626,WX9673,CRC_OUT_2_20);
  nand NAND2_6169(II31627,WX9673,II31626);
  nand NAND2_6170(II31628,CRC_OUT_2_20,II31626);
  nand NAND2_6171(WX10296,II31627,II31628);
  nand NAND2_6172(II31633,WX9674,CRC_OUT_2_19);
  nand NAND2_6173(II31634,WX9674,II31633);
  nand NAND2_6174(II31635,CRC_OUT_2_19,II31633);
  nand NAND2_6175(WX10297,II31634,II31635);
  nand NAND2_6176(II31640,WX9675,CRC_OUT_2_18);
  nand NAND2_6177(II31641,WX9675,II31640);
  nand NAND2_6178(II31642,CRC_OUT_2_18,II31640);
  nand NAND2_6179(WX10298,II31641,II31642);
  nand NAND2_6180(II31647,WX9676,CRC_OUT_2_17);
  nand NAND2_6181(II31648,WX9676,II31647);
  nand NAND2_6182(II31649,CRC_OUT_2_17,II31647);
  nand NAND2_6183(WX10299,II31648,II31649);
  nand NAND2_6184(II31654,WX9677,CRC_OUT_2_16);
  nand NAND2_6185(II31655,WX9677,II31654);
  nand NAND2_6186(II31656,CRC_OUT_2_16,II31654);
  nand NAND2_6187(WX10300,II31655,II31656);
  nand NAND2_6188(II31661,WX9679,CRC_OUT_2_14);
  nand NAND2_6189(II31662,WX9679,II31661);
  nand NAND2_6190(II31663,CRC_OUT_2_14,II31661);
  nand NAND2_6191(WX10301,II31662,II31663);
  nand NAND2_6192(II31668,WX9680,CRC_OUT_2_13);
  nand NAND2_6193(II31669,WX9680,II31668);
  nand NAND2_6194(II31670,CRC_OUT_2_13,II31668);
  nand NAND2_6195(WX10302,II31669,II31670);
  nand NAND2_6196(II31675,WX9681,CRC_OUT_2_12);
  nand NAND2_6197(II31676,WX9681,II31675);
  nand NAND2_6198(II31677,CRC_OUT_2_12,II31675);
  nand NAND2_6199(WX10303,II31676,II31677);
  nand NAND2_6200(II31682,WX9682,CRC_OUT_2_11);
  nand NAND2_6201(II31683,WX9682,II31682);
  nand NAND2_6202(II31684,CRC_OUT_2_11,II31682);
  nand NAND2_6203(WX10304,II31683,II31684);
  nand NAND2_6204(II31689,WX9684,CRC_OUT_2_9);
  nand NAND2_6205(II31690,WX9684,II31689);
  nand NAND2_6206(II31691,CRC_OUT_2_9,II31689);
  nand NAND2_6207(WX10305,II31690,II31691);
  nand NAND2_6208(II31696,WX9685,CRC_OUT_2_8);
  nand NAND2_6209(II31697,WX9685,II31696);
  nand NAND2_6210(II31698,CRC_OUT_2_8,II31696);
  nand NAND2_6211(WX10306,II31697,II31698);
  nand NAND2_6212(II31703,WX9686,CRC_OUT_2_7);
  nand NAND2_6213(II31704,WX9686,II31703);
  nand NAND2_6214(II31705,CRC_OUT_2_7,II31703);
  nand NAND2_6215(WX10307,II31704,II31705);
  nand NAND2_6216(II31710,WX9687,CRC_OUT_2_6);
  nand NAND2_6217(II31711,WX9687,II31710);
  nand NAND2_6218(II31712,CRC_OUT_2_6,II31710);
  nand NAND2_6219(WX10308,II31711,II31712);
  nand NAND2_6220(II31717,WX9688,CRC_OUT_2_5);
  nand NAND2_6221(II31718,WX9688,II31717);
  nand NAND2_6222(II31719,CRC_OUT_2_5,II31717);
  nand NAND2_6223(WX10309,II31718,II31719);
  nand NAND2_6224(II31724,WX9689,CRC_OUT_2_4);
  nand NAND2_6225(II31725,WX9689,II31724);
  nand NAND2_6226(II31726,CRC_OUT_2_4,II31724);
  nand NAND2_6227(WX10310,II31725,II31726);
  nand NAND2_6228(II31731,WX9691,CRC_OUT_2_2);
  nand NAND2_6229(II31732,WX9691,II31731);
  nand NAND2_6230(II31733,CRC_OUT_2_2,II31731);
  nand NAND2_6231(WX10311,II31732,II31733);
  nand NAND2_6232(II31738,WX9692,CRC_OUT_2_1);
  nand NAND2_6233(II31739,WX9692,II31738);
  nand NAND2_6234(II31740,CRC_OUT_2_1,II31738);
  nand NAND2_6235(WX10312,II31739,II31740);
  nand NAND2_6236(II31745,WX9693,CRC_OUT_2_0);
  nand NAND2_6237(II31746,WX9693,II31745);
  nand NAND2_6238(II31747,CRC_OUT_2_0,II31745);
  nand NAND2_6239(WX10313,II31746,II31747);
  nand NAND2_6240(II34028,WX11345,WX10989);
  nand NAND2_6241(II34029,WX11345,II34028);
  nand NAND2_6242(II34030,WX10989,II34028);
  nand NAND2_6243(II34027,II34029,II34030);
  nand NAND2_6244(II34035,WX11053,II34027);
  nand NAND2_6245(II34036,WX11053,II34035);
  nand NAND2_6246(II34037,II34027,II34035);
  nand NAND2_6247(II34026,II34036,II34037);
  nand NAND2_6248(II34043,WX11117,WX11181);
  nand NAND2_6249(II34044,WX11117,II34043);
  nand NAND2_6250(II34045,WX11181,II34043);
  nand NAND2_6251(II34042,II34044,II34045);
  nand NAND2_6252(II34050,II34026,II34042);
  nand NAND2_6253(II34051,II34026,II34050);
  nand NAND2_6254(II34052,II34042,II34050);
  nand NAND2_6255(WX11244,II34051,II34052);
  nand NAND2_6256(II34059,WX11345,WX10991);
  nand NAND2_6257(II34060,WX11345,II34059);
  nand NAND2_6258(II34061,WX10991,II34059);
  nand NAND2_6259(II34058,II34060,II34061);
  nand NAND2_6260(II34066,WX11055,II34058);
  nand NAND2_6261(II34067,WX11055,II34066);
  nand NAND2_6262(II34068,II34058,II34066);
  nand NAND2_6263(II34057,II34067,II34068);
  nand NAND2_6264(II34074,WX11119,WX11183);
  nand NAND2_6265(II34075,WX11119,II34074);
  nand NAND2_6266(II34076,WX11183,II34074);
  nand NAND2_6267(II34073,II34075,II34076);
  nand NAND2_6268(II34081,II34057,II34073);
  nand NAND2_6269(II34082,II34057,II34081);
  nand NAND2_6270(II34083,II34073,II34081);
  nand NAND2_6271(WX11245,II34082,II34083);
  nand NAND2_6272(II34090,WX11345,WX10993);
  nand NAND2_6273(II34091,WX11345,II34090);
  nand NAND2_6274(II34092,WX10993,II34090);
  nand NAND2_6275(II34089,II34091,II34092);
  nand NAND2_6276(II34097,WX11057,II34089);
  nand NAND2_6277(II34098,WX11057,II34097);
  nand NAND2_6278(II34099,II34089,II34097);
  nand NAND2_6279(II34088,II34098,II34099);
  nand NAND2_6280(II34105,WX11121,WX11185);
  nand NAND2_6281(II34106,WX11121,II34105);
  nand NAND2_6282(II34107,WX11185,II34105);
  nand NAND2_6283(II34104,II34106,II34107);
  nand NAND2_6284(II34112,II34088,II34104);
  nand NAND2_6285(II34113,II34088,II34112);
  nand NAND2_6286(II34114,II34104,II34112);
  nand NAND2_6287(WX11246,II34113,II34114);
  nand NAND2_6288(II34121,WX11345,WX10995);
  nand NAND2_6289(II34122,WX11345,II34121);
  nand NAND2_6290(II34123,WX10995,II34121);
  nand NAND2_6291(II34120,II34122,II34123);
  nand NAND2_6292(II34128,WX11059,II34120);
  nand NAND2_6293(II34129,WX11059,II34128);
  nand NAND2_6294(II34130,II34120,II34128);
  nand NAND2_6295(II34119,II34129,II34130);
  nand NAND2_6296(II34136,WX11123,WX11187);
  nand NAND2_6297(II34137,WX11123,II34136);
  nand NAND2_6298(II34138,WX11187,II34136);
  nand NAND2_6299(II34135,II34137,II34138);
  nand NAND2_6300(II34143,II34119,II34135);
  nand NAND2_6301(II34144,II34119,II34143);
  nand NAND2_6302(II34145,II34135,II34143);
  nand NAND2_6303(WX11247,II34144,II34145);
  nand NAND2_6304(II34152,WX11345,WX10997);
  nand NAND2_6305(II34153,WX11345,II34152);
  nand NAND2_6306(II34154,WX10997,II34152);
  nand NAND2_6307(II34151,II34153,II34154);
  nand NAND2_6308(II34159,WX11061,II34151);
  nand NAND2_6309(II34160,WX11061,II34159);
  nand NAND2_6310(II34161,II34151,II34159);
  nand NAND2_6311(II34150,II34160,II34161);
  nand NAND2_6312(II34167,WX11125,WX11189);
  nand NAND2_6313(II34168,WX11125,II34167);
  nand NAND2_6314(II34169,WX11189,II34167);
  nand NAND2_6315(II34166,II34168,II34169);
  nand NAND2_6316(II34174,II34150,II34166);
  nand NAND2_6317(II34175,II34150,II34174);
  nand NAND2_6318(II34176,II34166,II34174);
  nand NAND2_6319(WX11248,II34175,II34176);
  nand NAND2_6320(II34183,WX11345,WX10999);
  nand NAND2_6321(II34184,WX11345,II34183);
  nand NAND2_6322(II34185,WX10999,II34183);
  nand NAND2_6323(II34182,II34184,II34185);
  nand NAND2_6324(II34190,WX11063,II34182);
  nand NAND2_6325(II34191,WX11063,II34190);
  nand NAND2_6326(II34192,II34182,II34190);
  nand NAND2_6327(II34181,II34191,II34192);
  nand NAND2_6328(II34198,WX11127,WX11191);
  nand NAND2_6329(II34199,WX11127,II34198);
  nand NAND2_6330(II34200,WX11191,II34198);
  nand NAND2_6331(II34197,II34199,II34200);
  nand NAND2_6332(II34205,II34181,II34197);
  nand NAND2_6333(II34206,II34181,II34205);
  nand NAND2_6334(II34207,II34197,II34205);
  nand NAND2_6335(WX11249,II34206,II34207);
  nand NAND2_6336(II34214,WX11345,WX11001);
  nand NAND2_6337(II34215,WX11345,II34214);
  nand NAND2_6338(II34216,WX11001,II34214);
  nand NAND2_6339(II34213,II34215,II34216);
  nand NAND2_6340(II34221,WX11065,II34213);
  nand NAND2_6341(II34222,WX11065,II34221);
  nand NAND2_6342(II34223,II34213,II34221);
  nand NAND2_6343(II34212,II34222,II34223);
  nand NAND2_6344(II34229,WX11129,WX11193);
  nand NAND2_6345(II34230,WX11129,II34229);
  nand NAND2_6346(II34231,WX11193,II34229);
  nand NAND2_6347(II34228,II34230,II34231);
  nand NAND2_6348(II34236,II34212,II34228);
  nand NAND2_6349(II34237,II34212,II34236);
  nand NAND2_6350(II34238,II34228,II34236);
  nand NAND2_6351(WX11250,II34237,II34238);
  nand NAND2_6352(II34245,WX11345,WX11003);
  nand NAND2_6353(II34246,WX11345,II34245);
  nand NAND2_6354(II34247,WX11003,II34245);
  nand NAND2_6355(II34244,II34246,II34247);
  nand NAND2_6356(II34252,WX11067,II34244);
  nand NAND2_6357(II34253,WX11067,II34252);
  nand NAND2_6358(II34254,II34244,II34252);
  nand NAND2_6359(II34243,II34253,II34254);
  nand NAND2_6360(II34260,WX11131,WX11195);
  nand NAND2_6361(II34261,WX11131,II34260);
  nand NAND2_6362(II34262,WX11195,II34260);
  nand NAND2_6363(II34259,II34261,II34262);
  nand NAND2_6364(II34267,II34243,II34259);
  nand NAND2_6365(II34268,II34243,II34267);
  nand NAND2_6366(II34269,II34259,II34267);
  nand NAND2_6367(WX11251,II34268,II34269);
  nand NAND2_6368(II34276,WX11345,WX11005);
  nand NAND2_6369(II34277,WX11345,II34276);
  nand NAND2_6370(II34278,WX11005,II34276);
  nand NAND2_6371(II34275,II34277,II34278);
  nand NAND2_6372(II34283,WX11069,II34275);
  nand NAND2_6373(II34284,WX11069,II34283);
  nand NAND2_6374(II34285,II34275,II34283);
  nand NAND2_6375(II34274,II34284,II34285);
  nand NAND2_6376(II34291,WX11133,WX11197);
  nand NAND2_6377(II34292,WX11133,II34291);
  nand NAND2_6378(II34293,WX11197,II34291);
  nand NAND2_6379(II34290,II34292,II34293);
  nand NAND2_6380(II34298,II34274,II34290);
  nand NAND2_6381(II34299,II34274,II34298);
  nand NAND2_6382(II34300,II34290,II34298);
  nand NAND2_6383(WX11252,II34299,II34300);
  nand NAND2_6384(II34307,WX11345,WX11007);
  nand NAND2_6385(II34308,WX11345,II34307);
  nand NAND2_6386(II34309,WX11007,II34307);
  nand NAND2_6387(II34306,II34308,II34309);
  nand NAND2_6388(II34314,WX11071,II34306);
  nand NAND2_6389(II34315,WX11071,II34314);
  nand NAND2_6390(II34316,II34306,II34314);
  nand NAND2_6391(II34305,II34315,II34316);
  nand NAND2_6392(II34322,WX11135,WX11199);
  nand NAND2_6393(II34323,WX11135,II34322);
  nand NAND2_6394(II34324,WX11199,II34322);
  nand NAND2_6395(II34321,II34323,II34324);
  nand NAND2_6396(II34329,II34305,II34321);
  nand NAND2_6397(II34330,II34305,II34329);
  nand NAND2_6398(II34331,II34321,II34329);
  nand NAND2_6399(WX11253,II34330,II34331);
  nand NAND2_6400(II34338,WX11345,WX11009);
  nand NAND2_6401(II34339,WX11345,II34338);
  nand NAND2_6402(II34340,WX11009,II34338);
  nand NAND2_6403(II34337,II34339,II34340);
  nand NAND2_6404(II34345,WX11073,II34337);
  nand NAND2_6405(II34346,WX11073,II34345);
  nand NAND2_6406(II34347,II34337,II34345);
  nand NAND2_6407(II34336,II34346,II34347);
  nand NAND2_6408(II34353,WX11137,WX11201);
  nand NAND2_6409(II34354,WX11137,II34353);
  nand NAND2_6410(II34355,WX11201,II34353);
  nand NAND2_6411(II34352,II34354,II34355);
  nand NAND2_6412(II34360,II34336,II34352);
  nand NAND2_6413(II34361,II34336,II34360);
  nand NAND2_6414(II34362,II34352,II34360);
  nand NAND2_6415(WX11254,II34361,II34362);
  nand NAND2_6416(II34369,WX11345,WX11011);
  nand NAND2_6417(II34370,WX11345,II34369);
  nand NAND2_6418(II34371,WX11011,II34369);
  nand NAND2_6419(II34368,II34370,II34371);
  nand NAND2_6420(II34376,WX11075,II34368);
  nand NAND2_6421(II34377,WX11075,II34376);
  nand NAND2_6422(II34378,II34368,II34376);
  nand NAND2_6423(II34367,II34377,II34378);
  nand NAND2_6424(II34384,WX11139,WX11203);
  nand NAND2_6425(II34385,WX11139,II34384);
  nand NAND2_6426(II34386,WX11203,II34384);
  nand NAND2_6427(II34383,II34385,II34386);
  nand NAND2_6428(II34391,II34367,II34383);
  nand NAND2_6429(II34392,II34367,II34391);
  nand NAND2_6430(II34393,II34383,II34391);
  nand NAND2_6431(WX11255,II34392,II34393);
  nand NAND2_6432(II34400,WX11345,WX11013);
  nand NAND2_6433(II34401,WX11345,II34400);
  nand NAND2_6434(II34402,WX11013,II34400);
  nand NAND2_6435(II34399,II34401,II34402);
  nand NAND2_6436(II34407,WX11077,II34399);
  nand NAND2_6437(II34408,WX11077,II34407);
  nand NAND2_6438(II34409,II34399,II34407);
  nand NAND2_6439(II34398,II34408,II34409);
  nand NAND2_6440(II34415,WX11141,WX11205);
  nand NAND2_6441(II34416,WX11141,II34415);
  nand NAND2_6442(II34417,WX11205,II34415);
  nand NAND2_6443(II34414,II34416,II34417);
  nand NAND2_6444(II34422,II34398,II34414);
  nand NAND2_6445(II34423,II34398,II34422);
  nand NAND2_6446(II34424,II34414,II34422);
  nand NAND2_6447(WX11256,II34423,II34424);
  nand NAND2_6448(II34431,WX11345,WX11015);
  nand NAND2_6449(II34432,WX11345,II34431);
  nand NAND2_6450(II34433,WX11015,II34431);
  nand NAND2_6451(II34430,II34432,II34433);
  nand NAND2_6452(II34438,WX11079,II34430);
  nand NAND2_6453(II34439,WX11079,II34438);
  nand NAND2_6454(II34440,II34430,II34438);
  nand NAND2_6455(II34429,II34439,II34440);
  nand NAND2_6456(II34446,WX11143,WX11207);
  nand NAND2_6457(II34447,WX11143,II34446);
  nand NAND2_6458(II34448,WX11207,II34446);
  nand NAND2_6459(II34445,II34447,II34448);
  nand NAND2_6460(II34453,II34429,II34445);
  nand NAND2_6461(II34454,II34429,II34453);
  nand NAND2_6462(II34455,II34445,II34453);
  nand NAND2_6463(WX11257,II34454,II34455);
  nand NAND2_6464(II34462,WX11345,WX11017);
  nand NAND2_6465(II34463,WX11345,II34462);
  nand NAND2_6466(II34464,WX11017,II34462);
  nand NAND2_6467(II34461,II34463,II34464);
  nand NAND2_6468(II34469,WX11081,II34461);
  nand NAND2_6469(II34470,WX11081,II34469);
  nand NAND2_6470(II34471,II34461,II34469);
  nand NAND2_6471(II34460,II34470,II34471);
  nand NAND2_6472(II34477,WX11145,WX11209);
  nand NAND2_6473(II34478,WX11145,II34477);
  nand NAND2_6474(II34479,WX11209,II34477);
  nand NAND2_6475(II34476,II34478,II34479);
  nand NAND2_6476(II34484,II34460,II34476);
  nand NAND2_6477(II34485,II34460,II34484);
  nand NAND2_6478(II34486,II34476,II34484);
  nand NAND2_6479(WX11258,II34485,II34486);
  nand NAND2_6480(II34493,WX11345,WX11019);
  nand NAND2_6481(II34494,WX11345,II34493);
  nand NAND2_6482(II34495,WX11019,II34493);
  nand NAND2_6483(II34492,II34494,II34495);
  nand NAND2_6484(II34500,WX11083,II34492);
  nand NAND2_6485(II34501,WX11083,II34500);
  nand NAND2_6486(II34502,II34492,II34500);
  nand NAND2_6487(II34491,II34501,II34502);
  nand NAND2_6488(II34508,WX11147,WX11211);
  nand NAND2_6489(II34509,WX11147,II34508);
  nand NAND2_6490(II34510,WX11211,II34508);
  nand NAND2_6491(II34507,II34509,II34510);
  nand NAND2_6492(II34515,II34491,II34507);
  nand NAND2_6493(II34516,II34491,II34515);
  nand NAND2_6494(II34517,II34507,II34515);
  nand NAND2_6495(WX11259,II34516,II34517);
  nand NAND2_6496(II34524,WX11346,WX11021);
  nand NAND2_6497(II34525,WX11346,II34524);
  nand NAND2_6498(II34526,WX11021,II34524);
  nand NAND2_6499(II34523,II34525,II34526);
  nand NAND2_6500(II34531,WX11085,II34523);
  nand NAND2_6501(II34532,WX11085,II34531);
  nand NAND2_6502(II34533,II34523,II34531);
  nand NAND2_6503(II34522,II34532,II34533);
  nand NAND2_6504(II34539,WX11149,WX11213);
  nand NAND2_6505(II34540,WX11149,II34539);
  nand NAND2_6506(II34541,WX11213,II34539);
  nand NAND2_6507(II34538,II34540,II34541);
  nand NAND2_6508(II34546,II34522,II34538);
  nand NAND2_6509(II34547,II34522,II34546);
  nand NAND2_6510(II34548,II34538,II34546);
  nand NAND2_6511(WX11260,II34547,II34548);
  nand NAND2_6512(II34555,WX11346,WX11023);
  nand NAND2_6513(II34556,WX11346,II34555);
  nand NAND2_6514(II34557,WX11023,II34555);
  nand NAND2_6515(II34554,II34556,II34557);
  nand NAND2_6516(II34562,WX11087,II34554);
  nand NAND2_6517(II34563,WX11087,II34562);
  nand NAND2_6518(II34564,II34554,II34562);
  nand NAND2_6519(II34553,II34563,II34564);
  nand NAND2_6520(II34570,WX11151,WX11215);
  nand NAND2_6521(II34571,WX11151,II34570);
  nand NAND2_6522(II34572,WX11215,II34570);
  nand NAND2_6523(II34569,II34571,II34572);
  nand NAND2_6524(II34577,II34553,II34569);
  nand NAND2_6525(II34578,II34553,II34577);
  nand NAND2_6526(II34579,II34569,II34577);
  nand NAND2_6527(WX11261,II34578,II34579);
  nand NAND2_6528(II34586,WX11346,WX11025);
  nand NAND2_6529(II34587,WX11346,II34586);
  nand NAND2_6530(II34588,WX11025,II34586);
  nand NAND2_6531(II34585,II34587,II34588);
  nand NAND2_6532(II34593,WX11089,II34585);
  nand NAND2_6533(II34594,WX11089,II34593);
  nand NAND2_6534(II34595,II34585,II34593);
  nand NAND2_6535(II34584,II34594,II34595);
  nand NAND2_6536(II34601,WX11153,WX11217);
  nand NAND2_6537(II34602,WX11153,II34601);
  nand NAND2_6538(II34603,WX11217,II34601);
  nand NAND2_6539(II34600,II34602,II34603);
  nand NAND2_6540(II34608,II34584,II34600);
  nand NAND2_6541(II34609,II34584,II34608);
  nand NAND2_6542(II34610,II34600,II34608);
  nand NAND2_6543(WX11262,II34609,II34610);
  nand NAND2_6544(II34617,WX11346,WX11027);
  nand NAND2_6545(II34618,WX11346,II34617);
  nand NAND2_6546(II34619,WX11027,II34617);
  nand NAND2_6547(II34616,II34618,II34619);
  nand NAND2_6548(II34624,WX11091,II34616);
  nand NAND2_6549(II34625,WX11091,II34624);
  nand NAND2_6550(II34626,II34616,II34624);
  nand NAND2_6551(II34615,II34625,II34626);
  nand NAND2_6552(II34632,WX11155,WX11219);
  nand NAND2_6553(II34633,WX11155,II34632);
  nand NAND2_6554(II34634,WX11219,II34632);
  nand NAND2_6555(II34631,II34633,II34634);
  nand NAND2_6556(II34639,II34615,II34631);
  nand NAND2_6557(II34640,II34615,II34639);
  nand NAND2_6558(II34641,II34631,II34639);
  nand NAND2_6559(WX11263,II34640,II34641);
  nand NAND2_6560(II34648,WX11346,WX11029);
  nand NAND2_6561(II34649,WX11346,II34648);
  nand NAND2_6562(II34650,WX11029,II34648);
  nand NAND2_6563(II34647,II34649,II34650);
  nand NAND2_6564(II34655,WX11093,II34647);
  nand NAND2_6565(II34656,WX11093,II34655);
  nand NAND2_6566(II34657,II34647,II34655);
  nand NAND2_6567(II34646,II34656,II34657);
  nand NAND2_6568(II34663,WX11157,WX11221);
  nand NAND2_6569(II34664,WX11157,II34663);
  nand NAND2_6570(II34665,WX11221,II34663);
  nand NAND2_6571(II34662,II34664,II34665);
  nand NAND2_6572(II34670,II34646,II34662);
  nand NAND2_6573(II34671,II34646,II34670);
  nand NAND2_6574(II34672,II34662,II34670);
  nand NAND2_6575(WX11264,II34671,II34672);
  nand NAND2_6576(II34679,WX11346,WX11031);
  nand NAND2_6577(II34680,WX11346,II34679);
  nand NAND2_6578(II34681,WX11031,II34679);
  nand NAND2_6579(II34678,II34680,II34681);
  nand NAND2_6580(II34686,WX11095,II34678);
  nand NAND2_6581(II34687,WX11095,II34686);
  nand NAND2_6582(II34688,II34678,II34686);
  nand NAND2_6583(II34677,II34687,II34688);
  nand NAND2_6584(II34694,WX11159,WX11223);
  nand NAND2_6585(II34695,WX11159,II34694);
  nand NAND2_6586(II34696,WX11223,II34694);
  nand NAND2_6587(II34693,II34695,II34696);
  nand NAND2_6588(II34701,II34677,II34693);
  nand NAND2_6589(II34702,II34677,II34701);
  nand NAND2_6590(II34703,II34693,II34701);
  nand NAND2_6591(WX11265,II34702,II34703);
  nand NAND2_6592(II34710,WX11346,WX11033);
  nand NAND2_6593(II34711,WX11346,II34710);
  nand NAND2_6594(II34712,WX11033,II34710);
  nand NAND2_6595(II34709,II34711,II34712);
  nand NAND2_6596(II34717,WX11097,II34709);
  nand NAND2_6597(II34718,WX11097,II34717);
  nand NAND2_6598(II34719,II34709,II34717);
  nand NAND2_6599(II34708,II34718,II34719);
  nand NAND2_6600(II34725,WX11161,WX11225);
  nand NAND2_6601(II34726,WX11161,II34725);
  nand NAND2_6602(II34727,WX11225,II34725);
  nand NAND2_6603(II34724,II34726,II34727);
  nand NAND2_6604(II34732,II34708,II34724);
  nand NAND2_6605(II34733,II34708,II34732);
  nand NAND2_6606(II34734,II34724,II34732);
  nand NAND2_6607(WX11266,II34733,II34734);
  nand NAND2_6608(II34741,WX11346,WX11035);
  nand NAND2_6609(II34742,WX11346,II34741);
  nand NAND2_6610(II34743,WX11035,II34741);
  nand NAND2_6611(II34740,II34742,II34743);
  nand NAND2_6612(II34748,WX11099,II34740);
  nand NAND2_6613(II34749,WX11099,II34748);
  nand NAND2_6614(II34750,II34740,II34748);
  nand NAND2_6615(II34739,II34749,II34750);
  nand NAND2_6616(II34756,WX11163,WX11227);
  nand NAND2_6617(II34757,WX11163,II34756);
  nand NAND2_6618(II34758,WX11227,II34756);
  nand NAND2_6619(II34755,II34757,II34758);
  nand NAND2_6620(II34763,II34739,II34755);
  nand NAND2_6621(II34764,II34739,II34763);
  nand NAND2_6622(II34765,II34755,II34763);
  nand NAND2_6623(WX11267,II34764,II34765);
  nand NAND2_6624(II34772,WX11346,WX11037);
  nand NAND2_6625(II34773,WX11346,II34772);
  nand NAND2_6626(II34774,WX11037,II34772);
  nand NAND2_6627(II34771,II34773,II34774);
  nand NAND2_6628(II34779,WX11101,II34771);
  nand NAND2_6629(II34780,WX11101,II34779);
  nand NAND2_6630(II34781,II34771,II34779);
  nand NAND2_6631(II34770,II34780,II34781);
  nand NAND2_6632(II34787,WX11165,WX11229);
  nand NAND2_6633(II34788,WX11165,II34787);
  nand NAND2_6634(II34789,WX11229,II34787);
  nand NAND2_6635(II34786,II34788,II34789);
  nand NAND2_6636(II34794,II34770,II34786);
  nand NAND2_6637(II34795,II34770,II34794);
  nand NAND2_6638(II34796,II34786,II34794);
  nand NAND2_6639(WX11268,II34795,II34796);
  nand NAND2_6640(II34803,WX11346,WX11039);
  nand NAND2_6641(II34804,WX11346,II34803);
  nand NAND2_6642(II34805,WX11039,II34803);
  nand NAND2_6643(II34802,II34804,II34805);
  nand NAND2_6644(II34810,WX11103,II34802);
  nand NAND2_6645(II34811,WX11103,II34810);
  nand NAND2_6646(II34812,II34802,II34810);
  nand NAND2_6647(II34801,II34811,II34812);
  nand NAND2_6648(II34818,WX11167,WX11231);
  nand NAND2_6649(II34819,WX11167,II34818);
  nand NAND2_6650(II34820,WX11231,II34818);
  nand NAND2_6651(II34817,II34819,II34820);
  nand NAND2_6652(II34825,II34801,II34817);
  nand NAND2_6653(II34826,II34801,II34825);
  nand NAND2_6654(II34827,II34817,II34825);
  nand NAND2_6655(WX11269,II34826,II34827);
  nand NAND2_6656(II34834,WX11346,WX11041);
  nand NAND2_6657(II34835,WX11346,II34834);
  nand NAND2_6658(II34836,WX11041,II34834);
  nand NAND2_6659(II34833,II34835,II34836);
  nand NAND2_6660(II34841,WX11105,II34833);
  nand NAND2_6661(II34842,WX11105,II34841);
  nand NAND2_6662(II34843,II34833,II34841);
  nand NAND2_6663(II34832,II34842,II34843);
  nand NAND2_6664(II34849,WX11169,WX11233);
  nand NAND2_6665(II34850,WX11169,II34849);
  nand NAND2_6666(II34851,WX11233,II34849);
  nand NAND2_6667(II34848,II34850,II34851);
  nand NAND2_6668(II34856,II34832,II34848);
  nand NAND2_6669(II34857,II34832,II34856);
  nand NAND2_6670(II34858,II34848,II34856);
  nand NAND2_6671(WX11270,II34857,II34858);
  nand NAND2_6672(II34865,WX11346,WX11043);
  nand NAND2_6673(II34866,WX11346,II34865);
  nand NAND2_6674(II34867,WX11043,II34865);
  nand NAND2_6675(II34864,II34866,II34867);
  nand NAND2_6676(II34872,WX11107,II34864);
  nand NAND2_6677(II34873,WX11107,II34872);
  nand NAND2_6678(II34874,II34864,II34872);
  nand NAND2_6679(II34863,II34873,II34874);
  nand NAND2_6680(II34880,WX11171,WX11235);
  nand NAND2_6681(II34881,WX11171,II34880);
  nand NAND2_6682(II34882,WX11235,II34880);
  nand NAND2_6683(II34879,II34881,II34882);
  nand NAND2_6684(II34887,II34863,II34879);
  nand NAND2_6685(II34888,II34863,II34887);
  nand NAND2_6686(II34889,II34879,II34887);
  nand NAND2_6687(WX11271,II34888,II34889);
  nand NAND2_6688(II34896,WX11346,WX11045);
  nand NAND2_6689(II34897,WX11346,II34896);
  nand NAND2_6690(II34898,WX11045,II34896);
  nand NAND2_6691(II34895,II34897,II34898);
  nand NAND2_6692(II34903,WX11109,II34895);
  nand NAND2_6693(II34904,WX11109,II34903);
  nand NAND2_6694(II34905,II34895,II34903);
  nand NAND2_6695(II34894,II34904,II34905);
  nand NAND2_6696(II34911,WX11173,WX11237);
  nand NAND2_6697(II34912,WX11173,II34911);
  nand NAND2_6698(II34913,WX11237,II34911);
  nand NAND2_6699(II34910,II34912,II34913);
  nand NAND2_6700(II34918,II34894,II34910);
  nand NAND2_6701(II34919,II34894,II34918);
  nand NAND2_6702(II34920,II34910,II34918);
  nand NAND2_6703(WX11272,II34919,II34920);
  nand NAND2_6704(II34927,WX11346,WX11047);
  nand NAND2_6705(II34928,WX11346,II34927);
  nand NAND2_6706(II34929,WX11047,II34927);
  nand NAND2_6707(II34926,II34928,II34929);
  nand NAND2_6708(II34934,WX11111,II34926);
  nand NAND2_6709(II34935,WX11111,II34934);
  nand NAND2_6710(II34936,II34926,II34934);
  nand NAND2_6711(II34925,II34935,II34936);
  nand NAND2_6712(II34942,WX11175,WX11239);
  nand NAND2_6713(II34943,WX11175,II34942);
  nand NAND2_6714(II34944,WX11239,II34942);
  nand NAND2_6715(II34941,II34943,II34944);
  nand NAND2_6716(II34949,II34925,II34941);
  nand NAND2_6717(II34950,II34925,II34949);
  nand NAND2_6718(II34951,II34941,II34949);
  nand NAND2_6719(WX11273,II34950,II34951);
  nand NAND2_6720(II34958,WX11346,WX11049);
  nand NAND2_6721(II34959,WX11346,II34958);
  nand NAND2_6722(II34960,WX11049,II34958);
  nand NAND2_6723(II34957,II34959,II34960);
  nand NAND2_6724(II34965,WX11113,II34957);
  nand NAND2_6725(II34966,WX11113,II34965);
  nand NAND2_6726(II34967,II34957,II34965);
  nand NAND2_6727(II34956,II34966,II34967);
  nand NAND2_6728(II34973,WX11177,WX11241);
  nand NAND2_6729(II34974,WX11177,II34973);
  nand NAND2_6730(II34975,WX11241,II34973);
  nand NAND2_6731(II34972,II34974,II34975);
  nand NAND2_6732(II34980,II34956,II34972);
  nand NAND2_6733(II34981,II34956,II34980);
  nand NAND2_6734(II34982,II34972,II34980);
  nand NAND2_6735(WX11274,II34981,II34982);
  nand NAND2_6736(II34989,WX11346,WX11051);
  nand NAND2_6737(II34990,WX11346,II34989);
  nand NAND2_6738(II34991,WX11051,II34989);
  nand NAND2_6739(II34988,II34990,II34991);
  nand NAND2_6740(II34996,WX11115,II34988);
  nand NAND2_6741(II34997,WX11115,II34996);
  nand NAND2_6742(II34998,II34988,II34996);
  nand NAND2_6743(II34987,II34997,II34998);
  nand NAND2_6744(II35004,WX11179,WX11243);
  nand NAND2_6745(II35005,WX11179,II35004);
  nand NAND2_6746(II35006,WX11243,II35004);
  nand NAND2_6747(II35003,II35005,II35006);
  nand NAND2_6748(II35011,II34987,II35003);
  nand NAND2_6749(II35012,II34987,II35011);
  nand NAND2_6750(II35013,II35003,II35011);
  nand NAND2_6751(WX11275,II35012,II35013);
  nand NAND2_6752(II35092,WX10924,WX10829);
  nand NAND2_6753(II35093,WX10924,II35092);
  nand NAND2_6754(II35094,WX10829,II35092);
  nand NAND2_6755(WX11350,II35093,II35094);
  nand NAND2_6756(II35105,WX10925,WX10831);
  nand NAND2_6757(II35106,WX10925,II35105);
  nand NAND2_6758(II35107,WX10831,II35105);
  nand NAND2_6759(WX11357,II35106,II35107);
  nand NAND2_6760(II35118,WX10926,WX10833);
  nand NAND2_6761(II35119,WX10926,II35118);
  nand NAND2_6762(II35120,WX10833,II35118);
  nand NAND2_6763(WX11364,II35119,II35120);
  nand NAND2_6764(II35131,WX10927,WX10835);
  nand NAND2_6765(II35132,WX10927,II35131);
  nand NAND2_6766(II35133,WX10835,II35131);
  nand NAND2_6767(WX11371,II35132,II35133);
  nand NAND2_6768(II35144,WX10928,WX10837);
  nand NAND2_6769(II35145,WX10928,II35144);
  nand NAND2_6770(II35146,WX10837,II35144);
  nand NAND2_6771(WX11378,II35145,II35146);
  nand NAND2_6772(II35157,WX10929,WX10839);
  nand NAND2_6773(II35158,WX10929,II35157);
  nand NAND2_6774(II35159,WX10839,II35157);
  nand NAND2_6775(WX11385,II35158,II35159);
  nand NAND2_6776(II35170,WX10930,WX10841);
  nand NAND2_6777(II35171,WX10930,II35170);
  nand NAND2_6778(II35172,WX10841,II35170);
  nand NAND2_6779(WX11392,II35171,II35172);
  nand NAND2_6780(II35183,WX10931,WX10843);
  nand NAND2_6781(II35184,WX10931,II35183);
  nand NAND2_6782(II35185,WX10843,II35183);
  nand NAND2_6783(WX11399,II35184,II35185);
  nand NAND2_6784(II35196,WX10932,WX10845);
  nand NAND2_6785(II35197,WX10932,II35196);
  nand NAND2_6786(II35198,WX10845,II35196);
  nand NAND2_6787(WX11406,II35197,II35198);
  nand NAND2_6788(II35209,WX10933,WX10847);
  nand NAND2_6789(II35210,WX10933,II35209);
  nand NAND2_6790(II35211,WX10847,II35209);
  nand NAND2_6791(WX11413,II35210,II35211);
  nand NAND2_6792(II35222,WX10934,WX10849);
  nand NAND2_6793(II35223,WX10934,II35222);
  nand NAND2_6794(II35224,WX10849,II35222);
  nand NAND2_6795(WX11420,II35223,II35224);
  nand NAND2_6796(II35235,WX10935,WX10851);
  nand NAND2_6797(II35236,WX10935,II35235);
  nand NAND2_6798(II35237,WX10851,II35235);
  nand NAND2_6799(WX11427,II35236,II35237);
  nand NAND2_6800(II35248,WX10936,WX10853);
  nand NAND2_6801(II35249,WX10936,II35248);
  nand NAND2_6802(II35250,WX10853,II35248);
  nand NAND2_6803(WX11434,II35249,II35250);
  nand NAND2_6804(II35261,WX10937,WX10855);
  nand NAND2_6805(II35262,WX10937,II35261);
  nand NAND2_6806(II35263,WX10855,II35261);
  nand NAND2_6807(WX11441,II35262,II35263);
  nand NAND2_6808(II35274,WX10938,WX10857);
  nand NAND2_6809(II35275,WX10938,II35274);
  nand NAND2_6810(II35276,WX10857,II35274);
  nand NAND2_6811(WX11448,II35275,II35276);
  nand NAND2_6812(II35287,WX10939,WX10859);
  nand NAND2_6813(II35288,WX10939,II35287);
  nand NAND2_6814(II35289,WX10859,II35287);
  nand NAND2_6815(WX11455,II35288,II35289);
  nand NAND2_6816(II35300,WX10940,WX10861);
  nand NAND2_6817(II35301,WX10940,II35300);
  nand NAND2_6818(II35302,WX10861,II35300);
  nand NAND2_6819(WX11462,II35301,II35302);
  nand NAND2_6820(II35313,WX10941,WX10863);
  nand NAND2_6821(II35314,WX10941,II35313);
  nand NAND2_6822(II35315,WX10863,II35313);
  nand NAND2_6823(WX11469,II35314,II35315);
  nand NAND2_6824(II35326,WX10942,WX10865);
  nand NAND2_6825(II35327,WX10942,II35326);
  nand NAND2_6826(II35328,WX10865,II35326);
  nand NAND2_6827(WX11476,II35327,II35328);
  nand NAND2_6828(II35339,WX10943,WX10867);
  nand NAND2_6829(II35340,WX10943,II35339);
  nand NAND2_6830(II35341,WX10867,II35339);
  nand NAND2_6831(WX11483,II35340,II35341);
  nand NAND2_6832(II35352,WX10944,WX10869);
  nand NAND2_6833(II35353,WX10944,II35352);
  nand NAND2_6834(II35354,WX10869,II35352);
  nand NAND2_6835(WX11490,II35353,II35354);
  nand NAND2_6836(II35365,WX10945,WX10871);
  nand NAND2_6837(II35366,WX10945,II35365);
  nand NAND2_6838(II35367,WX10871,II35365);
  nand NAND2_6839(WX11497,II35366,II35367);
  nand NAND2_6840(II35378,WX10946,WX10873);
  nand NAND2_6841(II35379,WX10946,II35378);
  nand NAND2_6842(II35380,WX10873,II35378);
  nand NAND2_6843(WX11504,II35379,II35380);
  nand NAND2_6844(II35391,WX10947,WX10875);
  nand NAND2_6845(II35392,WX10947,II35391);
  nand NAND2_6846(II35393,WX10875,II35391);
  nand NAND2_6847(WX11511,II35392,II35393);
  nand NAND2_6848(II35404,WX10948,WX10877);
  nand NAND2_6849(II35405,WX10948,II35404);
  nand NAND2_6850(II35406,WX10877,II35404);
  nand NAND2_6851(WX11518,II35405,II35406);
  nand NAND2_6852(II35417,WX10949,WX10879);
  nand NAND2_6853(II35418,WX10949,II35417);
  nand NAND2_6854(II35419,WX10879,II35417);
  nand NAND2_6855(WX11525,II35418,II35419);
  nand NAND2_6856(II35430,WX10950,WX10881);
  nand NAND2_6857(II35431,WX10950,II35430);
  nand NAND2_6858(II35432,WX10881,II35430);
  nand NAND2_6859(WX11532,II35431,II35432);
  nand NAND2_6860(II35443,WX10951,WX10883);
  nand NAND2_6861(II35444,WX10951,II35443);
  nand NAND2_6862(II35445,WX10883,II35443);
  nand NAND2_6863(WX11539,II35444,II35445);
  nand NAND2_6864(II35456,WX10952,WX10885);
  nand NAND2_6865(II35457,WX10952,II35456);
  nand NAND2_6866(II35458,WX10885,II35456);
  nand NAND2_6867(WX11546,II35457,II35458);
  nand NAND2_6868(II35469,WX10953,WX10887);
  nand NAND2_6869(II35470,WX10953,II35469);
  nand NAND2_6870(II35471,WX10887,II35469);
  nand NAND2_6871(WX11553,II35470,II35471);
  nand NAND2_6872(II35482,WX10954,WX10889);
  nand NAND2_6873(II35483,WX10954,II35482);
  nand NAND2_6874(II35484,WX10889,II35482);
  nand NAND2_6875(WX11560,II35483,II35484);
  nand NAND2_6876(II35495,WX10955,WX10891);
  nand NAND2_6877(II35496,WX10955,II35495);
  nand NAND2_6878(II35497,WX10891,II35495);
  nand NAND2_6879(WX11567,II35496,II35497);
  nand NAND2_6880(II35510,WX10971,CRC_OUT_1_31);
  nand NAND2_6881(II35511,WX10971,II35510);
  nand NAND2_6882(II35512,CRC_OUT_1_31,II35510);
  nand NAND2_6883(II35509,II35511,II35512);
  nand NAND2_6884(II35517,CRC_OUT_1_15,II35509);
  nand NAND2_6885(II35518,CRC_OUT_1_15,II35517);
  nand NAND2_6886(II35519,II35509,II35517);
  nand NAND2_6887(WX11575,II35518,II35519);
  nand NAND2_6888(II35525,WX10976,CRC_OUT_1_31);
  nand NAND2_6889(II35526,WX10976,II35525);
  nand NAND2_6890(II35527,CRC_OUT_1_31,II35525);
  nand NAND2_6891(II35524,II35526,II35527);
  nand NAND2_6892(II35532,CRC_OUT_1_10,II35524);
  nand NAND2_6893(II35533,CRC_OUT_1_10,II35532);
  nand NAND2_6894(II35534,II35524,II35532);
  nand NAND2_6895(WX11576,II35533,II35534);
  nand NAND2_6896(II35540,WX10983,CRC_OUT_1_31);
  nand NAND2_6897(II35541,WX10983,II35540);
  nand NAND2_6898(II35542,CRC_OUT_1_31,II35540);
  nand NAND2_6899(II35539,II35541,II35542);
  nand NAND2_6900(II35547,CRC_OUT_1_3,II35539);
  nand NAND2_6901(II35548,CRC_OUT_1_3,II35547);
  nand NAND2_6902(II35549,II35539,II35547);
  nand NAND2_6903(WX11577,II35548,II35549);
  nand NAND2_6904(II35554,WX10987,CRC_OUT_1_31);
  nand NAND2_6905(II35555,WX10987,II35554);
  nand NAND2_6906(II35556,CRC_OUT_1_31,II35554);
  nand NAND2_6907(WX11578,II35555,II35556);
  nand NAND2_6908(II35561,WX10956,CRC_OUT_1_30);
  nand NAND2_6909(II35562,WX10956,II35561);
  nand NAND2_6910(II35563,CRC_OUT_1_30,II35561);
  nand NAND2_6911(WX11579,II35562,II35563);
  nand NAND2_6912(II35568,WX10957,CRC_OUT_1_29);
  nand NAND2_6913(II35569,WX10957,II35568);
  nand NAND2_6914(II35570,CRC_OUT_1_29,II35568);
  nand NAND2_6915(WX11580,II35569,II35570);
  nand NAND2_6916(II35575,WX10958,CRC_OUT_1_28);
  nand NAND2_6917(II35576,WX10958,II35575);
  nand NAND2_6918(II35577,CRC_OUT_1_28,II35575);
  nand NAND2_6919(WX11581,II35576,II35577);
  nand NAND2_6920(II35582,WX10959,CRC_OUT_1_27);
  nand NAND2_6921(II35583,WX10959,II35582);
  nand NAND2_6922(II35584,CRC_OUT_1_27,II35582);
  nand NAND2_6923(WX11582,II35583,II35584);
  nand NAND2_6924(II35589,WX10960,CRC_OUT_1_26);
  nand NAND2_6925(II35590,WX10960,II35589);
  nand NAND2_6926(II35591,CRC_OUT_1_26,II35589);
  nand NAND2_6927(WX11583,II35590,II35591);
  nand NAND2_6928(II35596,WX10961,CRC_OUT_1_25);
  nand NAND2_6929(II35597,WX10961,II35596);
  nand NAND2_6930(II35598,CRC_OUT_1_25,II35596);
  nand NAND2_6931(WX11584,II35597,II35598);
  nand NAND2_6932(II35603,WX10962,CRC_OUT_1_24);
  nand NAND2_6933(II35604,WX10962,II35603);
  nand NAND2_6934(II35605,CRC_OUT_1_24,II35603);
  nand NAND2_6935(WX11585,II35604,II35605);
  nand NAND2_6936(II35610,WX10963,CRC_OUT_1_23);
  nand NAND2_6937(II35611,WX10963,II35610);
  nand NAND2_6938(II35612,CRC_OUT_1_23,II35610);
  nand NAND2_6939(WX11586,II35611,II35612);
  nand NAND2_6940(II35617,WX10964,CRC_OUT_1_22);
  nand NAND2_6941(II35618,WX10964,II35617);
  nand NAND2_6942(II35619,CRC_OUT_1_22,II35617);
  nand NAND2_6943(WX11587,II35618,II35619);
  nand NAND2_6944(II35624,WX10965,CRC_OUT_1_21);
  nand NAND2_6945(II35625,WX10965,II35624);
  nand NAND2_6946(II35626,CRC_OUT_1_21,II35624);
  nand NAND2_6947(WX11588,II35625,II35626);
  nand NAND2_6948(II35631,WX10966,CRC_OUT_1_20);
  nand NAND2_6949(II35632,WX10966,II35631);
  nand NAND2_6950(II35633,CRC_OUT_1_20,II35631);
  nand NAND2_6951(WX11589,II35632,II35633);
  nand NAND2_6952(II35638,WX10967,CRC_OUT_1_19);
  nand NAND2_6953(II35639,WX10967,II35638);
  nand NAND2_6954(II35640,CRC_OUT_1_19,II35638);
  nand NAND2_6955(WX11590,II35639,II35640);
  nand NAND2_6956(II35645,WX10968,CRC_OUT_1_18);
  nand NAND2_6957(II35646,WX10968,II35645);
  nand NAND2_6958(II35647,CRC_OUT_1_18,II35645);
  nand NAND2_6959(WX11591,II35646,II35647);
  nand NAND2_6960(II35652,WX10969,CRC_OUT_1_17);
  nand NAND2_6961(II35653,WX10969,II35652);
  nand NAND2_6962(II35654,CRC_OUT_1_17,II35652);
  nand NAND2_6963(WX11592,II35653,II35654);
  nand NAND2_6964(II35659,WX10970,CRC_OUT_1_16);
  nand NAND2_6965(II35660,WX10970,II35659);
  nand NAND2_6966(II35661,CRC_OUT_1_16,II35659);
  nand NAND2_6967(WX11593,II35660,II35661);
  nand NAND2_6968(II35666,WX10972,CRC_OUT_1_14);
  nand NAND2_6969(II35667,WX10972,II35666);
  nand NAND2_6970(II35668,CRC_OUT_1_14,II35666);
  nand NAND2_6971(WX11594,II35667,II35668);
  nand NAND2_6972(II35673,WX10973,CRC_OUT_1_13);
  nand NAND2_6973(II35674,WX10973,II35673);
  nand NAND2_6974(II35675,CRC_OUT_1_13,II35673);
  nand NAND2_6975(WX11595,II35674,II35675);
  nand NAND2_6976(II35680,WX10974,CRC_OUT_1_12);
  nand NAND2_6977(II35681,WX10974,II35680);
  nand NAND2_6978(II35682,CRC_OUT_1_12,II35680);
  nand NAND2_6979(WX11596,II35681,II35682);
  nand NAND2_6980(II35687,WX10975,CRC_OUT_1_11);
  nand NAND2_6981(II35688,WX10975,II35687);
  nand NAND2_6982(II35689,CRC_OUT_1_11,II35687);
  nand NAND2_6983(WX11597,II35688,II35689);
  nand NAND2_6984(II35694,WX10977,CRC_OUT_1_9);
  nand NAND2_6985(II35695,WX10977,II35694);
  nand NAND2_6986(II35696,CRC_OUT_1_9,II35694);
  nand NAND2_6987(WX11598,II35695,II35696);
  nand NAND2_6988(II35701,WX10978,CRC_OUT_1_8);
  nand NAND2_6989(II35702,WX10978,II35701);
  nand NAND2_6990(II35703,CRC_OUT_1_8,II35701);
  nand NAND2_6991(WX11599,II35702,II35703);
  nand NAND2_6992(II35708,WX10979,CRC_OUT_1_7);
  nand NAND2_6993(II35709,WX10979,II35708);
  nand NAND2_6994(II35710,CRC_OUT_1_7,II35708);
  nand NAND2_6995(WX11600,II35709,II35710);
  nand NAND2_6996(II35715,WX10980,CRC_OUT_1_6);
  nand NAND2_6997(II35716,WX10980,II35715);
  nand NAND2_6998(II35717,CRC_OUT_1_6,II35715);
  nand NAND2_6999(WX11601,II35716,II35717);
  nand NAND2_7000(II35722,WX10981,CRC_OUT_1_5);
  nand NAND2_7001(II35723,WX10981,II35722);
  nand NAND2_7002(II35724,CRC_OUT_1_5,II35722);
  nand NAND2_7003(WX11602,II35723,II35724);
  nand NAND2_7004(II35729,WX10982,CRC_OUT_1_4);
  nand NAND2_7005(II35730,WX10982,II35729);
  nand NAND2_7006(II35731,CRC_OUT_1_4,II35729);
  nand NAND2_7007(WX11603,II35730,II35731);
  nand NAND2_7008(II35736,WX10984,CRC_OUT_1_2);
  nand NAND2_7009(II35737,WX10984,II35736);
  nand NAND2_7010(II35738,CRC_OUT_1_2,II35736);
  nand NAND2_7011(WX11604,II35737,II35738);
  nand NAND2_7012(II35743,WX10985,CRC_OUT_1_1);
  nand NAND2_7013(II35744,WX10985,II35743);
  nand NAND2_7014(II35745,CRC_OUT_1_1,II35743);
  nand NAND2_7015(WX11605,II35744,II35745);
  nand NAND2_7016(II35750,WX10986,CRC_OUT_1_0);
  nand NAND2_7017(II35751,WX10986,II35750);
  nand NAND2_7018(II35752,CRC_OUT_1_0,II35750);
  nand NAND2_7019(WX11606,II35751,II35752);

endmodule//# 35 inputs
//# 320 outputs
//# 1728 D-type flipflops
//# 3861 inverters
//# 12204 gates (4032 ANDs + 7020 NANDs + 1152 ORs + 0 NORs)

module dff (CK,Q,D);
input CK,D;
output Q;

  wire NM,NCK;
  trireg NQ,M;

  nmos N7 (M,D,NCK);
  not P3 (NM,M);
  nmos N9 (NQ,NM,CK);
  not P5 (Q,NQ);
  not P1 (NCK,CK);

endmodule

module s35932(GND,VDD,CK,CRC_OUT_1_0,CRC_OUT_1_1,CRC_OUT_1_10,CRC_OUT_1_11,
  CRC_OUT_1_12,CRC_OUT_1_13,CRC_OUT_1_14,CRC_OUT_1_15,CRC_OUT_1_16,CRC_OUT_1_17,
  CRC_OUT_1_18,CRC_OUT_1_19,CRC_OUT_1_2,CRC_OUT_1_20,CRC_OUT_1_21,CRC_OUT_1_22,
  CRC_OUT_1_23,CRC_OUT_1_24,CRC_OUT_1_25,CRC_OUT_1_26,CRC_OUT_1_27,
  CRC_OUT_1_28,CRC_OUT_1_29,CRC_OUT_1_3,CRC_OUT_1_30,CRC_OUT_1_31,CRC_OUT_1_4,
  CRC_OUT_1_5,CRC_OUT_1_6,CRC_OUT_1_7,CRC_OUT_1_8,CRC_OUT_1_9,CRC_OUT_2_0,
  CRC_OUT_2_1,CRC_OUT_2_10,CRC_OUT_2_11,CRC_OUT_2_12,CRC_OUT_2_13,CRC_OUT_2_14,
  CRC_OUT_2_15,CRC_OUT_2_16,CRC_OUT_2_17,CRC_OUT_2_18,CRC_OUT_2_19,CRC_OUT_2_2,
  CRC_OUT_2_20,CRC_OUT_2_21,CRC_OUT_2_22,CRC_OUT_2_23,CRC_OUT_2_24,
  CRC_OUT_2_25,CRC_OUT_2_26,CRC_OUT_2_27,CRC_OUT_2_28,CRC_OUT_2_29,CRC_OUT_2_3,
  CRC_OUT_2_30,CRC_OUT_2_31,CRC_OUT_2_4,CRC_OUT_2_5,CRC_OUT_2_6,CRC_OUT_2_7,
  CRC_OUT_2_8,CRC_OUT_2_9,CRC_OUT_3_0,CRC_OUT_3_1,CRC_OUT_3_10,CRC_OUT_3_11,
  CRC_OUT_3_12,CRC_OUT_3_13,CRC_OUT_3_14,CRC_OUT_3_15,CRC_OUT_3_16,
  CRC_OUT_3_17,CRC_OUT_3_18,CRC_OUT_3_19,CRC_OUT_3_2,CRC_OUT_3_20,CRC_OUT_3_21,
  CRC_OUT_3_22,CRC_OUT_3_23,CRC_OUT_3_24,CRC_OUT_3_25,CRC_OUT_3_26,
  CRC_OUT_3_27,CRC_OUT_3_28,CRC_OUT_3_29,CRC_OUT_3_3,CRC_OUT_3_30,CRC_OUT_3_31,
  CRC_OUT_3_4,CRC_OUT_3_5,CRC_OUT_3_6,CRC_OUT_3_7,CRC_OUT_3_8,CRC_OUT_3_9,
  CRC_OUT_4_0,CRC_OUT_4_1,CRC_OUT_4_10,CRC_OUT_4_11,CRC_OUT_4_12,CRC_OUT_4_13,
  CRC_OUT_4_14,CRC_OUT_4_15,CRC_OUT_4_16,CRC_OUT_4_17,CRC_OUT_4_18,
  CRC_OUT_4_19,CRC_OUT_4_2,CRC_OUT_4_20,CRC_OUT_4_21,CRC_OUT_4_22,CRC_OUT_4_23,
  CRC_OUT_4_24,CRC_OUT_4_25,CRC_OUT_4_26,CRC_OUT_4_27,CRC_OUT_4_28,
  CRC_OUT_4_29,CRC_OUT_4_3,CRC_OUT_4_30,CRC_OUT_4_31,CRC_OUT_4_4,CRC_OUT_4_5,
  CRC_OUT_4_6,CRC_OUT_4_7,CRC_OUT_4_8,CRC_OUT_4_9,CRC_OUT_5_0,CRC_OUT_5_1,
  CRC_OUT_5_10,CRC_OUT_5_11,CRC_OUT_5_12,CRC_OUT_5_13,CRC_OUT_5_14,
  CRC_OUT_5_15,CRC_OUT_5_16,CRC_OUT_5_17,CRC_OUT_5_18,CRC_OUT_5_19,CRC_OUT_5_2,
  CRC_OUT_5_20,CRC_OUT_5_21,CRC_OUT_5_22,CRC_OUT_5_23,CRC_OUT_5_24,
  CRC_OUT_5_25,CRC_OUT_5_26,CRC_OUT_5_27,CRC_OUT_5_28,CRC_OUT_5_29,CRC_OUT_5_3,
  CRC_OUT_5_30,CRC_OUT_5_31,CRC_OUT_5_4,CRC_OUT_5_5,CRC_OUT_5_6,CRC_OUT_5_7,
  CRC_OUT_5_8,CRC_OUT_5_9,CRC_OUT_6_0,CRC_OUT_6_1,CRC_OUT_6_10,CRC_OUT_6_11,
  CRC_OUT_6_12,CRC_OUT_6_13,CRC_OUT_6_14,CRC_OUT_6_15,CRC_OUT_6_16,
  CRC_OUT_6_17,CRC_OUT_6_18,CRC_OUT_6_19,CRC_OUT_6_2,CRC_OUT_6_20,CRC_OUT_6_21,
  CRC_OUT_6_22,CRC_OUT_6_23,CRC_OUT_6_24,CRC_OUT_6_25,CRC_OUT_6_26,
  CRC_OUT_6_27,CRC_OUT_6_28,CRC_OUT_6_29,CRC_OUT_6_3,CRC_OUT_6_30,CRC_OUT_6_31,
  CRC_OUT_6_4,CRC_OUT_6_5,CRC_OUT_6_6,CRC_OUT_6_7,CRC_OUT_6_8,CRC_OUT_6_9,
  CRC_OUT_7_0,CRC_OUT_7_1,CRC_OUT_7_10,CRC_OUT_7_11,CRC_OUT_7_12,CRC_OUT_7_13,
  CRC_OUT_7_14,CRC_OUT_7_15,CRC_OUT_7_16,CRC_OUT_7_17,CRC_OUT_7_18,
  CRC_OUT_7_19,CRC_OUT_7_2,CRC_OUT_7_20,CRC_OUT_7_21,CRC_OUT_7_22,CRC_OUT_7_23,
  CRC_OUT_7_24,CRC_OUT_7_25,CRC_OUT_7_26,CRC_OUT_7_27,CRC_OUT_7_28,
  CRC_OUT_7_29,CRC_OUT_7_3,CRC_OUT_7_30,CRC_OUT_7_31,CRC_OUT_7_4,CRC_OUT_7_5,
  CRC_OUT_7_6,CRC_OUT_7_7,CRC_OUT_7_8,CRC_OUT_7_9,CRC_OUT_8_0,CRC_OUT_8_1,
  CRC_OUT_8_10,CRC_OUT_8_11,CRC_OUT_8_12,CRC_OUT_8_13,CRC_OUT_8_14,
  CRC_OUT_8_15,CRC_OUT_8_16,CRC_OUT_8_17,CRC_OUT_8_18,CRC_OUT_8_19,CRC_OUT_8_2,
  CRC_OUT_8_20,CRC_OUT_8_21,CRC_OUT_8_22,CRC_OUT_8_23,CRC_OUT_8_24,
  CRC_OUT_8_25,CRC_OUT_8_26,CRC_OUT_8_27,CRC_OUT_8_28,CRC_OUT_8_29,CRC_OUT_8_3,
  CRC_OUT_8_30,CRC_OUT_8_31,CRC_OUT_8_4,CRC_OUT_8_5,CRC_OUT_8_6,CRC_OUT_8_7,
  CRC_OUT_8_8,CRC_OUT_8_9,CRC_OUT_9_0,CRC_OUT_9_1,CRC_OUT_9_10,CRC_OUT_9_11,
  CRC_OUT_9_12,CRC_OUT_9_13,CRC_OUT_9_14,CRC_OUT_9_15,CRC_OUT_9_16,
  CRC_OUT_9_17,CRC_OUT_9_18,CRC_OUT_9_19,CRC_OUT_9_2,CRC_OUT_9_20,CRC_OUT_9_21,
  CRC_OUT_9_22,CRC_OUT_9_23,CRC_OUT_9_24,CRC_OUT_9_25,CRC_OUT_9_26,
  CRC_OUT_9_27,CRC_OUT_9_28,CRC_OUT_9_29,CRC_OUT_9_3,CRC_OUT_9_30,CRC_OUT_9_31,
  CRC_OUT_9_4,CRC_OUT_9_5,CRC_OUT_9_6,CRC_OUT_9_7,CRC_OUT_9_8,CRC_OUT_9_9,
  DATA_0_0,DATA_0_1,DATA_0_10,DATA_0_11,DATA_0_12,DATA_0_13,DATA_0_14,
  DATA_0_15,DATA_0_16,DATA_0_17,DATA_0_18,DATA_0_19,DATA_0_2,DATA_0_20,
  DATA_0_21,DATA_0_22,DATA_0_23,DATA_0_24,DATA_0_25,DATA_0_26,DATA_0_27,
  DATA_0_28,DATA_0_29,DATA_0_3,DATA_0_30,DATA_0_31,DATA_0_4,DATA_0_5,DATA_0_6,
  DATA_0_7,DATA_0_8,DATA_0_9,DATA_9_0,DATA_9_1,DATA_9_10,DATA_9_11,DATA_9_12,
  DATA_9_13,DATA_9_14,DATA_9_15,DATA_9_16,DATA_9_17,DATA_9_18,DATA_9_19,
  DATA_9_2,DATA_9_20,DATA_9_21,DATA_9_22,DATA_9_23,DATA_9_24,DATA_9_25,
  DATA_9_26,DATA_9_27,DATA_9_28,DATA_9_29,DATA_9_3,DATA_9_30,DATA_9_31,
  DATA_9_4,DATA_9_5,DATA_9_6,DATA_9_7,DATA_9_8,DATA_9_9,RESET,TM0,TM1);
input GND,VDD,CK,DATA_0_31,DATA_0_30,DATA_0_29,DATA_0_28,DATA_0_27,DATA_0_26,
  DATA_0_25,
  DATA_0_24,DATA_0_23,DATA_0_22,DATA_0_21,DATA_0_20,DATA_0_19,DATA_0_18,
  DATA_0_17,DATA_0_16,DATA_0_15,DATA_0_14,DATA_0_13,DATA_0_12,DATA_0_11,
  DATA_0_10,DATA_0_9,DATA_0_8,DATA_0_7,DATA_0_6,DATA_0_5,DATA_0_4,DATA_0_3,
  DATA_0_2,DATA_0_1,DATA_0_0,RESET,TM1,TM0;
output DATA_9_31,DATA_9_30,DATA_9_29,DATA_9_28,DATA_9_27,DATA_9_26,DATA_9_25,
  DATA_9_24,DATA_9_23,DATA_9_22,DATA_9_21,DATA_9_20,DATA_9_19,DATA_9_18,
  DATA_9_17,DATA_9_16,DATA_9_15,DATA_9_14,DATA_9_13,DATA_9_12,DATA_9_11,
  DATA_9_10,DATA_9_9,DATA_9_8,DATA_9_7,DATA_9_6,DATA_9_5,DATA_9_4,DATA_9_3,
  DATA_9_2,DATA_9_1,DATA_9_0,CRC_OUT_9_0,CRC_OUT_9_1,CRC_OUT_9_2,CRC_OUT_9_3,
  CRC_OUT_9_4,CRC_OUT_9_5,CRC_OUT_9_6,CRC_OUT_9_7,CRC_OUT_9_8,CRC_OUT_9_9,
  CRC_OUT_9_10,CRC_OUT_9_11,CRC_OUT_9_12,CRC_OUT_9_13,CRC_OUT_9_14,
  CRC_OUT_9_15,CRC_OUT_9_16,CRC_OUT_9_17,CRC_OUT_9_18,CRC_OUT_9_19,
  CRC_OUT_9_20,CRC_OUT_9_21,CRC_OUT_9_22,CRC_OUT_9_23,CRC_OUT_9_24,
  CRC_OUT_9_25,CRC_OUT_9_26,CRC_OUT_9_27,CRC_OUT_9_28,CRC_OUT_9_29,
  CRC_OUT_9_30,CRC_OUT_9_31,CRC_OUT_8_0,CRC_OUT_8_1,CRC_OUT_8_2,CRC_OUT_8_3,
  CRC_OUT_8_4,CRC_OUT_8_5,CRC_OUT_8_6,CRC_OUT_8_7,CRC_OUT_8_8,CRC_OUT_8_9,
  CRC_OUT_8_10,CRC_OUT_8_11,CRC_OUT_8_12,CRC_OUT_8_13,CRC_OUT_8_14,
  CRC_OUT_8_15,CRC_OUT_8_16,CRC_OUT_8_17,CRC_OUT_8_18,CRC_OUT_8_19,
  CRC_OUT_8_20,CRC_OUT_8_21,CRC_OUT_8_22,CRC_OUT_8_23,CRC_OUT_8_24,
  CRC_OUT_8_25,CRC_OUT_8_26,CRC_OUT_8_27,CRC_OUT_8_28,CRC_OUT_8_29,
  CRC_OUT_8_30,CRC_OUT_8_31,CRC_OUT_7_0,CRC_OUT_7_1,CRC_OUT_7_2,CRC_OUT_7_3,
  CRC_OUT_7_4,CRC_OUT_7_5,CRC_OUT_7_6,CRC_OUT_7_7,CRC_OUT_7_8,CRC_OUT_7_9,
  CRC_OUT_7_10,CRC_OUT_7_11,CRC_OUT_7_12,CRC_OUT_7_13,CRC_OUT_7_14,
  CRC_OUT_7_15,CRC_OUT_7_16,CRC_OUT_7_17,CRC_OUT_7_18,CRC_OUT_7_19,
  CRC_OUT_7_20,CRC_OUT_7_21,CRC_OUT_7_22,CRC_OUT_7_23,CRC_OUT_7_24,
  CRC_OUT_7_25,CRC_OUT_7_26,CRC_OUT_7_27,CRC_OUT_7_28,CRC_OUT_7_29,
  CRC_OUT_7_30,CRC_OUT_7_31,CRC_OUT_6_0,CRC_OUT_6_1,CRC_OUT_6_2,CRC_OUT_6_3,
  CRC_OUT_6_4,CRC_OUT_6_5,CRC_OUT_6_6,CRC_OUT_6_7,CRC_OUT_6_8,CRC_OUT_6_9,
  CRC_OUT_6_10,CRC_OUT_6_11,CRC_OUT_6_12,CRC_OUT_6_13,CRC_OUT_6_14,
  CRC_OUT_6_15,CRC_OUT_6_16,CRC_OUT_6_17,CRC_OUT_6_18,CRC_OUT_6_19,
  CRC_OUT_6_20,CRC_OUT_6_21,CRC_OUT_6_22,CRC_OUT_6_23,CRC_OUT_6_24,
  CRC_OUT_6_25,CRC_OUT_6_26,CRC_OUT_6_27,CRC_OUT_6_28,CRC_OUT_6_29,
  CRC_OUT_6_30,CRC_OUT_6_31,CRC_OUT_5_0,CRC_OUT_5_1,CRC_OUT_5_2,CRC_OUT_5_3,
  CRC_OUT_5_4,CRC_OUT_5_5,CRC_OUT_5_6,CRC_OUT_5_7,CRC_OUT_5_8,CRC_OUT_5_9,
  CRC_OUT_5_10,CRC_OUT_5_11,CRC_OUT_5_12,CRC_OUT_5_13,CRC_OUT_5_14,
  CRC_OUT_5_15,CRC_OUT_5_16,CRC_OUT_5_17,CRC_OUT_5_18,CRC_OUT_5_19,
  CRC_OUT_5_20,CRC_OUT_5_21,CRC_OUT_5_22,CRC_OUT_5_23,CRC_OUT_5_24,
  CRC_OUT_5_25,CRC_OUT_5_26,CRC_OUT_5_27,CRC_OUT_5_28,CRC_OUT_5_29,
  CRC_OUT_5_30,CRC_OUT_5_31,CRC_OUT_4_0,CRC_OUT_4_1,CRC_OUT_4_2,CRC_OUT_4_3,
  CRC_OUT_4_4,CRC_OUT_4_5,CRC_OUT_4_6,CRC_OUT_4_7,CRC_OUT_4_8,CRC_OUT_4_9,
  CRC_OUT_4_10,CRC_OUT_4_11,CRC_OUT_4_12,CRC_OUT_4_13,CRC_OUT_4_14,
  CRC_OUT_4_15,CRC_OUT_4_16,CRC_OUT_4_17,CRC_OUT_4_18,CRC_OUT_4_19,
  CRC_OUT_4_20,CRC_OUT_4_21,CRC_OUT_4_22,CRC_OUT_4_23,CRC_OUT_4_24,
  CRC_OUT_4_25,CRC_OUT_4_26,CRC_OUT_4_27,CRC_OUT_4_28,CRC_OUT_4_29,
  CRC_OUT_4_30,CRC_OUT_4_31,CRC_OUT_3_0,CRC_OUT_3_1,CRC_OUT_3_2,CRC_OUT_3_3,
  CRC_OUT_3_4,CRC_OUT_3_5,CRC_OUT_3_6,CRC_OUT_3_7,CRC_OUT_3_8,CRC_OUT_3_9,
  CRC_OUT_3_10,CRC_OUT_3_11,CRC_OUT_3_12,CRC_OUT_3_13,CRC_OUT_3_14,
  CRC_OUT_3_15,CRC_OUT_3_16,CRC_OUT_3_17,CRC_OUT_3_18,CRC_OUT_3_19,
  CRC_OUT_3_20,CRC_OUT_3_21,CRC_OUT_3_22,CRC_OUT_3_23,CRC_OUT_3_24,
  CRC_OUT_3_25,CRC_OUT_3_26,CRC_OUT_3_27,CRC_OUT_3_28,CRC_OUT_3_29,
  CRC_OUT_3_30,CRC_OUT_3_31,CRC_OUT_2_0,CRC_OUT_2_1,CRC_OUT_2_2,CRC_OUT_2_3,
  CRC_OUT_2_4,CRC_OUT_2_5,CRC_OUT_2_6,CRC_OUT_2_7,CRC_OUT_2_8,CRC_OUT_2_9,
  CRC_OUT_2_10,CRC_OUT_2_11,CRC_OUT_2_12,CRC_OUT_2_13,CRC_OUT_2_14,
  CRC_OUT_2_15,CRC_OUT_2_16,CRC_OUT_2_17,CRC_OUT_2_18,CRC_OUT_2_19,
  CRC_OUT_2_20,CRC_OUT_2_21,CRC_OUT_2_22,CRC_OUT_2_23,CRC_OUT_2_24,
  CRC_OUT_2_25,CRC_OUT_2_26,CRC_OUT_2_27,CRC_OUT_2_28,CRC_OUT_2_29,
  CRC_OUT_2_30,CRC_OUT_2_31,CRC_OUT_1_0,CRC_OUT_1_1,CRC_OUT_1_2,CRC_OUT_1_3,
  CRC_OUT_1_4,CRC_OUT_1_5,CRC_OUT_1_6,CRC_OUT_1_7,CRC_OUT_1_8,CRC_OUT_1_9,
  CRC_OUT_1_10,CRC_OUT_1_11,CRC_OUT_1_12,CRC_OUT_1_13,CRC_OUT_1_14,
  CRC_OUT_1_15,CRC_OUT_1_16,CRC_OUT_1_17,CRC_OUT_1_18,CRC_OUT_1_19,
  CRC_OUT_1_20,CRC_OUT_1_21,CRC_OUT_1_22,CRC_OUT_1_23,CRC_OUT_1_24,
  CRC_OUT_1_25,CRC_OUT_1_26,CRC_OUT_1_27,CRC_OUT_1_28,CRC_OUT_1_29,
  CRC_OUT_1_30,CRC_OUT_1_31;

  wire WX485,WX484,WX487,WX486,WX489,WX488,WX491,WX490,WX493,WX492,WX495,WX494,
    WX497,WX496,WX499,WX498,WX501,WX500,WX503,WX502,WX505,WX504,WX507,WX506,
    WX509,WX508,WX511,WX510,WX513,WX512,WX515,WX514,WX517,WX516,WX519,WX518,
    WX521,WX520,WX523,WX522,WX525,WX524,WX527,WX526,WX529,WX528,WX531,WX530,
    WX533,WX532,WX535,WX534,WX537,WX536,WX539,WX538,WX541,WX540,WX543,WX542,
    WX545,WX544,WX547,WX546,WX645,WX644,WX647,WX646,WX649,WX648,WX651,WX650,
    WX653,WX652,WX655,WX654,WX657,WX656,WX659,WX658,WX661,WX660,WX663,WX662,
    WX665,WX664,WX667,WX666,WX669,WX668,WX671,WX670,WX673,WX672,WX675,WX674,
    WX677,WX676,WX679,WX678,WX681,WX680,WX683,WX682,WX685,WX684,WX687,WX686,
    WX689,WX688,WX691,WX690,WX693,WX692,WX695,WX694,WX697,WX696,WX699,WX698,
    WX701,WX700,WX703,WX702,WX705,WX704,WX707,WX706,WX709,WX708,WX711,WX710,
    WX713,WX712,WX715,WX714,WX717,WX716,WX719,WX718,WX721,WX720,WX723,WX722,
    WX725,WX724,WX727,WX726,WX729,WX728,WX731,WX730,WX733,WX732,WX735,WX734,
    WX737,WX736,WX739,WX738,WX741,WX740,WX743,WX742,WX745,WX744,WX747,WX746,
    WX749,WX748,WX751,WX750,WX753,WX752,WX755,WX754,WX757,WX756,WX759,WX758,
    WX761,WX760,WX763,WX762,WX765,WX764,WX767,WX766,WX769,WX768,WX771,WX770,
    WX773,WX772,WX775,WX774,WX777,WX776,WX779,WX778,WX781,WX780,WX783,WX782,
    WX785,WX784,WX787,WX786,WX789,WX788,WX791,WX790,WX793,WX792,WX795,WX794,
    WX797,WX796,WX799,WX798,WX801,WX800,WX803,WX802,WX805,WX804,WX807,WX806,
    WX809,WX808,WX811,WX810,WX813,WX812,WX815,WX814,WX817,WX816,WX819,WX818,
    WX821,WX820,WX823,WX822,WX825,WX824,WX827,WX826,WX829,WX828,WX831,WX830,
    WX833,WX832,WX835,WX834,WX837,WX836,WX839,WX838,WX841,WX840,WX843,WX842,
    WX845,WX844,WX847,WX846,WX849,WX848,WX851,WX850,WX853,WX852,WX855,WX854,
    WX857,WX856,WX859,WX858,WX861,WX860,WX863,WX862,WX865,WX864,WX867,WX866,
    WX869,WX868,WX871,WX870,WX873,WX872,WX875,WX874,WX877,WX876,WX879,WX878,
    WX881,WX880,WX883,WX882,WX885,WX884,WX887,WX886,WX889,WX888,WX891,WX890,
    WX893,WX892,WX895,WX894,WX897,WX896,WX899,WX898,WX1264,WX1266,WX1268,
    WX1270,WX1272,WX1274,WX1276,WX1278,WX1280,WX1282,WX1284,WX1286,WX1288,
    WX1290,WX1292,WX1294,WX1296,WX1298,WX1300,WX1302,WX1304,WX1306,WX1308,
    WX1310,WX1312,WX1314,WX1316,WX1318,WX1320,WX1322,WX1324,WX1326,WX1778,
    WX1777,WX1780,WX1779,WX1782,WX1781,WX1784,WX1783,WX1786,WX1785,WX1788,
    WX1787,WX1790,WX1789,WX1792,WX1791,WX1794,WX1793,WX1796,WX1795,WX1798,
    WX1797,WX1800,WX1799,WX1802,WX1801,WX1804,WX1803,WX1806,WX1805,WX1808,
    WX1807,WX1810,WX1809,WX1812,WX1811,WX1814,WX1813,WX1816,WX1815,WX1818,
    WX1817,WX1820,WX1819,WX1822,WX1821,WX1824,WX1823,WX1826,WX1825,WX1828,
    WX1827,WX1830,WX1829,WX1832,WX1831,WX1834,WX1833,WX1836,WX1835,WX1838,
    WX1837,WX1840,WX1839,WX1938,WX1937,WX1940,WX1939,WX1942,WX1941,WX1944,
    WX1943,WX1946,WX1945,WX1948,WX1947,WX1950,WX1949,WX1952,WX1951,WX1954,
    WX1953,WX1956,WX1955,WX1958,WX1957,WX1960,WX1959,WX1962,WX1961,WX1964,
    WX1963,WX1966,WX1965,WX1968,WX1967,WX1970,WX1969,WX1972,WX1971,WX1974,
    WX1973,WX1976,WX1975,WX1978,WX1977,WX1980,WX1979,WX1982,WX1981,WX1984,
    WX1983,WX1986,WX1985,WX1988,WX1987,WX1990,WX1989,WX1992,WX1991,WX1994,
    WX1993,WX1996,WX1995,WX1998,WX1997,WX2000,WX1999,WX2002,WX2001,WX2004,
    WX2003,WX2006,WX2005,WX2008,WX2007,WX2010,WX2009,WX2012,WX2011,WX2014,
    WX2013,WX2016,WX2015,WX2018,WX2017,WX2020,WX2019,WX2022,WX2021,WX2024,
    WX2023,WX2026,WX2025,WX2028,WX2027,WX2030,WX2029,WX2032,WX2031,WX2034,
    WX2033,WX2036,WX2035,WX2038,WX2037,WX2040,WX2039,WX2042,WX2041,WX2044,
    WX2043,WX2046,WX2045,WX2048,WX2047,WX2050,WX2049,WX2052,WX2051,WX2054,
    WX2053,WX2056,WX2055,WX2058,WX2057,WX2060,WX2059,WX2062,WX2061,WX2064,
    WX2063,WX2066,WX2065,WX2068,WX2067,WX2070,WX2069,WX2072,WX2071,WX2074,
    WX2073,WX2076,WX2075,WX2078,WX2077,WX2080,WX2079,WX2082,WX2081,WX2084,
    WX2083,WX2086,WX2085,WX2088,WX2087,WX2090,WX2089,WX2092,WX2091,WX2094,
    WX2093,WX2096,WX2095,WX2098,WX2097,WX2100,WX2099,WX2102,WX2101,WX2104,
    WX2103,WX2106,WX2105,WX2108,WX2107,WX2110,WX2109,WX2112,WX2111,WX2114,
    WX2113,WX2116,WX2115,WX2118,WX2117,WX2120,WX2119,WX2122,WX2121,WX2124,
    WX2123,WX2126,WX2125,WX2128,WX2127,WX2130,WX2129,WX2132,WX2131,WX2134,
    WX2133,WX2136,WX2135,WX2138,WX2137,WX2140,WX2139,WX2142,WX2141,WX2144,
    WX2143,WX2146,WX2145,WX2148,WX2147,WX2150,WX2149,WX2152,WX2151,WX2154,
    WX2153,WX2156,WX2155,WX2158,WX2157,WX2160,WX2159,WX2162,WX2161,WX2164,
    WX2163,WX2166,WX2165,WX2168,WX2167,WX2170,WX2169,WX2172,WX2171,WX2174,
    WX2173,WX2176,WX2175,WX2178,WX2177,WX2180,WX2179,WX2182,WX2181,WX2184,
    WX2183,WX2186,WX2185,WX2188,WX2187,WX2190,WX2189,WX2192,WX2191,WX2557,
    WX2559,WX2561,WX2563,WX2565,WX2567,WX2569,WX2571,WX2573,WX2575,WX2577,
    WX2579,WX2581,WX2583,WX2585,WX2587,WX2589,WX2591,WX2593,WX2595,WX2597,
    WX2599,WX2601,WX2603,WX2605,WX2607,WX2609,WX2611,WX2613,WX2615,WX2617,
    WX2619,WX3071,WX3070,WX3073,WX3072,WX3075,WX3074,WX3077,WX3076,WX3079,
    WX3078,WX3081,WX3080,WX3083,WX3082,WX3085,WX3084,WX3087,WX3086,WX3089,
    WX3088,WX3091,WX3090,WX3093,WX3092,WX3095,WX3094,WX3097,WX3096,WX3099,
    WX3098,WX3101,WX3100,WX3103,WX3102,WX3105,WX3104,WX3107,WX3106,WX3109,
    WX3108,WX3111,WX3110,WX3113,WX3112,WX3115,WX3114,WX3117,WX3116,WX3119,
    WX3118,WX3121,WX3120,WX3123,WX3122,WX3125,WX3124,WX3127,WX3126,WX3129,
    WX3128,WX3131,WX3130,WX3133,WX3132,WX3231,WX3230,WX3233,WX3232,WX3235,
    WX3234,WX3237,WX3236,WX3239,WX3238,WX3241,WX3240,WX3243,WX3242,WX3245,
    WX3244,WX3247,WX3246,WX3249,WX3248,WX3251,WX3250,WX3253,WX3252,WX3255,
    WX3254,WX3257,WX3256,WX3259,WX3258,WX3261,WX3260,WX3263,WX3262,WX3265,
    WX3264,WX3267,WX3266,WX3269,WX3268,WX3271,WX3270,WX3273,WX3272,WX3275,
    WX3274,WX3277,WX3276,WX3279,WX3278,WX3281,WX3280,WX3283,WX3282,WX3285,
    WX3284,WX3287,WX3286,WX3289,WX3288,WX3291,WX3290,WX3293,WX3292,WX3295,
    WX3294,WX3297,WX3296,WX3299,WX3298,WX3301,WX3300,WX3303,WX3302,WX3305,
    WX3304,WX3307,WX3306,WX3309,WX3308,WX3311,WX3310,WX3313,WX3312,WX3315,
    WX3314,WX3317,WX3316,WX3319,WX3318,WX3321,WX3320,WX3323,WX3322,WX3325,
    WX3324,WX3327,WX3326,WX3329,WX3328,WX3331,WX3330,WX3333,WX3332,WX3335,
    WX3334,WX3337,WX3336,WX3339,WX3338,WX3341,WX3340,WX3343,WX3342,WX3345,
    WX3344,WX3347,WX3346,WX3349,WX3348,WX3351,WX3350,WX3353,WX3352,WX3355,
    WX3354,WX3357,WX3356,WX3359,WX3358,WX3361,WX3360,WX3363,WX3362,WX3365,
    WX3364,WX3367,WX3366,WX3369,WX3368,WX3371,WX3370,WX3373,WX3372,WX3375,
    WX3374,WX3377,WX3376,WX3379,WX3378,WX3381,WX3380,WX3383,WX3382,WX3385,
    WX3384,WX3387,WX3386,WX3389,WX3388,WX3391,WX3390,WX3393,WX3392,WX3395,
    WX3394,WX3397,WX3396,WX3399,WX3398,WX3401,WX3400,WX3403,WX3402,WX3405,
    WX3404,WX3407,WX3406,WX3409,WX3408,WX3411,WX3410,WX3413,WX3412,WX3415,
    WX3414,WX3417,WX3416,WX3419,WX3418,WX3421,WX3420,WX3423,WX3422,WX3425,
    WX3424,WX3427,WX3426,WX3429,WX3428,WX3431,WX3430,WX3433,WX3432,WX3435,
    WX3434,WX3437,WX3436,WX3439,WX3438,WX3441,WX3440,WX3443,WX3442,WX3445,
    WX3444,WX3447,WX3446,WX3449,WX3448,WX3451,WX3450,WX3453,WX3452,WX3455,
    WX3454,WX3457,WX3456,WX3459,WX3458,WX3461,WX3460,WX3463,WX3462,WX3465,
    WX3464,WX3467,WX3466,WX3469,WX3468,WX3471,WX3470,WX3473,WX3472,WX3475,
    WX3474,WX3477,WX3476,WX3479,WX3478,WX3481,WX3480,WX3483,WX3482,WX3485,
    WX3484,WX3850,WX3852,WX3854,WX3856,WX3858,WX3860,WX3862,WX3864,WX3866,
    WX3868,WX3870,WX3872,WX3874,WX3876,WX3878,WX3880,WX3882,WX3884,WX3886,
    WX3888,WX3890,WX3892,WX3894,WX3896,WX3898,WX3900,WX3902,WX3904,WX3906,
    WX3908,WX3910,WX3912,WX4364,WX4363,WX4366,WX4365,WX4368,WX4367,WX4370,
    WX4369,WX4372,WX4371,WX4374,WX4373,WX4376,WX4375,WX4378,WX4377,WX4380,
    WX4379,WX4382,WX4381,WX4384,WX4383,WX4386,WX4385,WX4388,WX4387,WX4390,
    WX4389,WX4392,WX4391,WX4394,WX4393,WX4396,WX4395,WX4398,WX4397,WX4400,
    WX4399,WX4402,WX4401,WX4404,WX4403,WX4406,WX4405,WX4408,WX4407,WX4410,
    WX4409,WX4412,WX4411,WX4414,WX4413,WX4416,WX4415,WX4418,WX4417,WX4420,
    WX4419,WX4422,WX4421,WX4424,WX4423,WX4426,WX4425,WX4524,WX4523,WX4526,
    WX4525,WX4528,WX4527,WX4530,WX4529,WX4532,WX4531,WX4534,WX4533,WX4536,
    WX4535,WX4538,WX4537,WX4540,WX4539,WX4542,WX4541,WX4544,WX4543,WX4546,
    WX4545,WX4548,WX4547,WX4550,WX4549,WX4552,WX4551,WX4554,WX4553,WX4556,
    WX4555,WX4558,WX4557,WX4560,WX4559,WX4562,WX4561,WX4564,WX4563,WX4566,
    WX4565,WX4568,WX4567,WX4570,WX4569,WX4572,WX4571,WX4574,WX4573,WX4576,
    WX4575,WX4578,WX4577,WX4580,WX4579,WX4582,WX4581,WX4584,WX4583,WX4586,
    WX4585,WX4588,WX4587,WX4590,WX4589,WX4592,WX4591,WX4594,WX4593,WX4596,
    WX4595,WX4598,WX4597,WX4600,WX4599,WX4602,WX4601,WX4604,WX4603,WX4606,
    WX4605,WX4608,WX4607,WX4610,WX4609,WX4612,WX4611,WX4614,WX4613,WX4616,
    WX4615,WX4618,WX4617,WX4620,WX4619,WX4622,WX4621,WX4624,WX4623,WX4626,
    WX4625,WX4628,WX4627,WX4630,WX4629,WX4632,WX4631,WX4634,WX4633,WX4636,
    WX4635,WX4638,WX4637,WX4640,WX4639,WX4642,WX4641,WX4644,WX4643,WX4646,
    WX4645,WX4648,WX4647,WX4650,WX4649,WX4652,WX4651,WX4654,WX4653,WX4656,
    WX4655,WX4658,WX4657,WX4660,WX4659,WX4662,WX4661,WX4664,WX4663,WX4666,
    WX4665,WX4668,WX4667,WX4670,WX4669,WX4672,WX4671,WX4674,WX4673,WX4676,
    WX4675,WX4678,WX4677,WX4680,WX4679,WX4682,WX4681,WX4684,WX4683,WX4686,
    WX4685,WX4688,WX4687,WX4690,WX4689,WX4692,WX4691,WX4694,WX4693,WX4696,
    WX4695,WX4698,WX4697,WX4700,WX4699,WX4702,WX4701,WX4704,WX4703,WX4706,
    WX4705,WX4708,WX4707,WX4710,WX4709,WX4712,WX4711,WX4714,WX4713,WX4716,
    WX4715,WX4718,WX4717,WX4720,WX4719,WX4722,WX4721,WX4724,WX4723,WX4726,
    WX4725,WX4728,WX4727,WX4730,WX4729,WX4732,WX4731,WX4734,WX4733,WX4736,
    WX4735,WX4738,WX4737,WX4740,WX4739,WX4742,WX4741,WX4744,WX4743,WX4746,
    WX4745,WX4748,WX4747,WX4750,WX4749,WX4752,WX4751,WX4754,WX4753,WX4756,
    WX4755,WX4758,WX4757,WX4760,WX4759,WX4762,WX4761,WX4764,WX4763,WX4766,
    WX4765,WX4768,WX4767,WX4770,WX4769,WX4772,WX4771,WX4774,WX4773,WX4776,
    WX4775,WX4778,WX4777,WX5143,WX5145,WX5147,WX5149,WX5151,WX5153,WX5155,
    WX5157,WX5159,WX5161,WX5163,WX5165,WX5167,WX5169,WX5171,WX5173,WX5175,
    WX5177,WX5179,WX5181,WX5183,WX5185,WX5187,WX5189,WX5191,WX5193,WX5195,
    WX5197,WX5199,WX5201,WX5203,WX5205,WX5657,WX5656,WX5659,WX5658,WX5661,
    WX5660,WX5663,WX5662,WX5665,WX5664,WX5667,WX5666,WX5669,WX5668,WX5671,
    WX5670,WX5673,WX5672,WX5675,WX5674,WX5677,WX5676,WX5679,WX5678,WX5681,
    WX5680,WX5683,WX5682,WX5685,WX5684,WX5687,WX5686,WX5689,WX5688,WX5691,
    WX5690,WX5693,WX5692,WX5695,WX5694,WX5697,WX5696,WX5699,WX5698,WX5701,
    WX5700,WX5703,WX5702,WX5705,WX5704,WX5707,WX5706,WX5709,WX5708,WX5711,
    WX5710,WX5713,WX5712,WX5715,WX5714,WX5717,WX5716,WX5719,WX5718,WX5817,
    WX5816,WX5819,WX5818,WX5821,WX5820,WX5823,WX5822,WX5825,WX5824,WX5827,
    WX5826,WX5829,WX5828,WX5831,WX5830,WX5833,WX5832,WX5835,WX5834,WX5837,
    WX5836,WX5839,WX5838,WX5841,WX5840,WX5843,WX5842,WX5845,WX5844,WX5847,
    WX5846,WX5849,WX5848,WX5851,WX5850,WX5853,WX5852,WX5855,WX5854,WX5857,
    WX5856,WX5859,WX5858,WX5861,WX5860,WX5863,WX5862,WX5865,WX5864,WX5867,
    WX5866,WX5869,WX5868,WX5871,WX5870,WX5873,WX5872,WX5875,WX5874,WX5877,
    WX5876,WX5879,WX5878,WX5881,WX5880,WX5883,WX5882,WX5885,WX5884,WX5887,
    WX5886,WX5889,WX5888,WX5891,WX5890,WX5893,WX5892,WX5895,WX5894,WX5897,
    WX5896,WX5899,WX5898,WX5901,WX5900,WX5903,WX5902,WX5905,WX5904,WX5907,
    WX5906,WX5909,WX5908,WX5911,WX5910,WX5913,WX5912,WX5915,WX5914,WX5917,
    WX5916,WX5919,WX5918,WX5921,WX5920,WX5923,WX5922,WX5925,WX5924,WX5927,
    WX5926,WX5929,WX5928,WX5931,WX5930,WX5933,WX5932,WX5935,WX5934,WX5937,
    WX5936,WX5939,WX5938,WX5941,WX5940,WX5943,WX5942,WX5945,WX5944,WX5947,
    WX5946,WX5949,WX5948,WX5951,WX5950,WX5953,WX5952,WX5955,WX5954,WX5957,
    WX5956,WX5959,WX5958,WX5961,WX5960,WX5963,WX5962,WX5965,WX5964,WX5967,
    WX5966,WX5969,WX5968,WX5971,WX5970,WX5973,WX5972,WX5975,WX5974,WX5977,
    WX5976,WX5979,WX5978,WX5981,WX5980,WX5983,WX5982,WX5985,WX5984,WX5987,
    WX5986,WX5989,WX5988,WX5991,WX5990,WX5993,WX5992,WX5995,WX5994,WX5997,
    WX5996,WX5999,WX5998,WX6001,WX6000,WX6003,WX6002,WX6005,WX6004,WX6007,
    WX6006,WX6009,WX6008,WX6011,WX6010,WX6013,WX6012,WX6015,WX6014,WX6017,
    WX6016,WX6019,WX6018,WX6021,WX6020,WX6023,WX6022,WX6025,WX6024,WX6027,
    WX6026,WX6029,WX6028,WX6031,WX6030,WX6033,WX6032,WX6035,WX6034,WX6037,
    WX6036,WX6039,WX6038,WX6041,WX6040,WX6043,WX6042,WX6045,WX6044,WX6047,
    WX6046,WX6049,WX6048,WX6051,WX6050,WX6053,WX6052,WX6055,WX6054,WX6057,
    WX6056,WX6059,WX6058,WX6061,WX6060,WX6063,WX6062,WX6065,WX6064,WX6067,
    WX6066,WX6069,WX6068,WX6071,WX6070,WX6436,WX6438,WX6440,WX6442,WX6444,
    WX6446,WX6448,WX6450,WX6452,WX6454,WX6456,WX6458,WX6460,WX6462,WX6464,
    WX6466,WX6468,WX6470,WX6472,WX6474,WX6476,WX6478,WX6480,WX6482,WX6484,
    WX6486,WX6488,WX6490,WX6492,WX6494,WX6496,WX6498,WX6950,WX6949,WX6952,
    WX6951,WX6954,WX6953,WX6956,WX6955,WX6958,WX6957,WX6960,WX6959,WX6962,
    WX6961,WX6964,WX6963,WX6966,WX6965,WX6968,WX6967,WX6970,WX6969,WX6972,
    WX6971,WX6974,WX6973,WX6976,WX6975,WX6978,WX6977,WX6980,WX6979,WX6982,
    WX6981,WX6984,WX6983,WX6986,WX6985,WX6988,WX6987,WX6990,WX6989,WX6992,
    WX6991,WX6994,WX6993,WX6996,WX6995,WX6998,WX6997,WX7000,WX6999,WX7002,
    WX7001,WX7004,WX7003,WX7006,WX7005,WX7008,WX7007,WX7010,WX7009,WX7012,
    WX7011,WX7110,WX7109,WX7112,WX7111,WX7114,WX7113,WX7116,WX7115,WX7118,
    WX7117,WX7120,WX7119,WX7122,WX7121,WX7124,WX7123,WX7126,WX7125,WX7128,
    WX7127,WX7130,WX7129,WX7132,WX7131,WX7134,WX7133,WX7136,WX7135,WX7138,
    WX7137,WX7140,WX7139,WX7142,WX7141,WX7144,WX7143,WX7146,WX7145,WX7148,
    WX7147,WX7150,WX7149,WX7152,WX7151,WX7154,WX7153,WX7156,WX7155,WX7158,
    WX7157,WX7160,WX7159,WX7162,WX7161,WX7164,WX7163,WX7166,WX7165,WX7168,
    WX7167,WX7170,WX7169,WX7172,WX7171,WX7174,WX7173,WX7176,WX7175,WX7178,
    WX7177,WX7180,WX7179,WX7182,WX7181,WX7184,WX7183,WX7186,WX7185,WX7188,
    WX7187,WX7190,WX7189,WX7192,WX7191,WX7194,WX7193,WX7196,WX7195,WX7198,
    WX7197,WX7200,WX7199,WX7202,WX7201,WX7204,WX7203,WX7206,WX7205,WX7208,
    WX7207,WX7210,WX7209,WX7212,WX7211,WX7214,WX7213,WX7216,WX7215,WX7218,
    WX7217,WX7220,WX7219,WX7222,WX7221,WX7224,WX7223,WX7226,WX7225,WX7228,
    WX7227,WX7230,WX7229,WX7232,WX7231,WX7234,WX7233,WX7236,WX7235,WX7238,
    WX7237,WX7240,WX7239,WX7242,WX7241,WX7244,WX7243,WX7246,WX7245,WX7248,
    WX7247,WX7250,WX7249,WX7252,WX7251,WX7254,WX7253,WX7256,WX7255,WX7258,
    WX7257,WX7260,WX7259,WX7262,WX7261,WX7264,WX7263,WX7266,WX7265,WX7268,
    WX7267,WX7270,WX7269,WX7272,WX7271,WX7274,WX7273,WX7276,WX7275,WX7278,
    WX7277,WX7280,WX7279,WX7282,WX7281,WX7284,WX7283,WX7286,WX7285,WX7288,
    WX7287,WX7290,WX7289,WX7292,WX7291,WX7294,WX7293,WX7296,WX7295,WX7298,
    WX7297,WX7300,WX7299,WX7302,WX7301,WX7304,WX7303,WX7306,WX7305,WX7308,
    WX7307,WX7310,WX7309,WX7312,WX7311,WX7314,WX7313,WX7316,WX7315,WX7318,
    WX7317,WX7320,WX7319,WX7322,WX7321,WX7324,WX7323,WX7326,WX7325,WX7328,
    WX7327,WX7330,WX7329,WX7332,WX7331,WX7334,WX7333,WX7336,WX7335,WX7338,
    WX7337,WX7340,WX7339,WX7342,WX7341,WX7344,WX7343,WX7346,WX7345,WX7348,
    WX7347,WX7350,WX7349,WX7352,WX7351,WX7354,WX7353,WX7356,WX7355,WX7358,
    WX7357,WX7360,WX7359,WX7362,WX7361,WX7364,WX7363,WX7729,WX7731,WX7733,
    WX7735,WX7737,WX7739,WX7741,WX7743,WX7745,WX7747,WX7749,WX7751,WX7753,
    WX7755,WX7757,WX7759,WX7761,WX7763,WX7765,WX7767,WX7769,WX7771,WX7773,
    WX7775,WX7777,WX7779,WX7781,WX7783,WX7785,WX7787,WX7789,WX7791,WX8243,
    WX8242,WX8245,WX8244,WX8247,WX8246,WX8249,WX8248,WX8251,WX8250,WX8253,
    WX8252,WX8255,WX8254,WX8257,WX8256,WX8259,WX8258,WX8261,WX8260,WX8263,
    WX8262,WX8265,WX8264,WX8267,WX8266,WX8269,WX8268,WX8271,WX8270,WX8273,
    WX8272,WX8275,WX8274,WX8277,WX8276,WX8279,WX8278,WX8281,WX8280,WX8283,
    WX8282,WX8285,WX8284,WX8287,WX8286,WX8289,WX8288,WX8291,WX8290,WX8293,
    WX8292,WX8295,WX8294,WX8297,WX8296,WX8299,WX8298,WX8301,WX8300,WX8303,
    WX8302,WX8305,WX8304,WX8403,WX8402,WX8405,WX8404,WX8407,WX8406,WX8409,
    WX8408,WX8411,WX8410,WX8413,WX8412,WX8415,WX8414,WX8417,WX8416,WX8419,
    WX8418,WX8421,WX8420,WX8423,WX8422,WX8425,WX8424,WX8427,WX8426,WX8429,
    WX8428,WX8431,WX8430,WX8433,WX8432,WX8435,WX8434,WX8437,WX8436,WX8439,
    WX8438,WX8441,WX8440,WX8443,WX8442,WX8445,WX8444,WX8447,WX8446,WX8449,
    WX8448,WX8451,WX8450,WX8453,WX8452,WX8455,WX8454,WX8457,WX8456,WX8459,
    WX8458,WX8461,WX8460,WX8463,WX8462,WX8465,WX8464,WX8467,WX8466,WX8469,
    WX8468,WX8471,WX8470,WX8473,WX8472,WX8475,WX8474,WX8477,WX8476,WX8479,
    WX8478,WX8481,WX8480,WX8483,WX8482,WX8485,WX8484,WX8487,WX8486,WX8489,
    WX8488,WX8491,WX8490,WX8493,WX8492,WX8495,WX8494,WX8497,WX8496,WX8499,
    WX8498,WX8501,WX8500,WX8503,WX8502,WX8505,WX8504,WX8507,WX8506,WX8509,
    WX8508,WX8511,WX8510,WX8513,WX8512,WX8515,WX8514,WX8517,WX8516,WX8519,
    WX8518,WX8521,WX8520,WX8523,WX8522,WX8525,WX8524,WX8527,WX8526,WX8529,
    WX8528,WX8531,WX8530,WX8533,WX8532,WX8535,WX8534,WX8537,WX8536,WX8539,
    WX8538,WX8541,WX8540,WX8543,WX8542,WX8545,WX8544,WX8547,WX8546,WX8549,
    WX8548,WX8551,WX8550,WX8553,WX8552,WX8555,WX8554,WX8557,WX8556,WX8559,
    WX8558,WX8561,WX8560,WX8563,WX8562,WX8565,WX8564,WX8567,WX8566,WX8569,
    WX8568,WX8571,WX8570,WX8573,WX8572,WX8575,WX8574,WX8577,WX8576,WX8579,
    WX8578,WX8581,WX8580,WX8583,WX8582,WX8585,WX8584,WX8587,WX8586,WX8589,
    WX8588,WX8591,WX8590,WX8593,WX8592,WX8595,WX8594,WX8597,WX8596,WX8599,
    WX8598,WX8601,WX8600,WX8603,WX8602,WX8605,WX8604,WX8607,WX8606,WX8609,
    WX8608,WX8611,WX8610,WX8613,WX8612,WX8615,WX8614,WX8617,WX8616,WX8619,
    WX8618,WX8621,WX8620,WX8623,WX8622,WX8625,WX8624,WX8627,WX8626,WX8629,
    WX8628,WX8631,WX8630,WX8633,WX8632,WX8635,WX8634,WX8637,WX8636,WX8639,
    WX8638,WX8641,WX8640,WX8643,WX8642,WX8645,WX8644,WX8647,WX8646,WX8649,
    WX8648,WX8651,WX8650,WX8653,WX8652,WX8655,WX8654,WX8657,WX8656,WX9022,
    WX9024,WX9026,WX9028,WX9030,WX9032,WX9034,WX9036,WX9038,WX9040,WX9042,
    WX9044,WX9046,WX9048,WX9050,WX9052,WX9054,WX9056,WX9058,WX9060,WX9062,
    WX9064,WX9066,WX9068,WX9070,WX9072,WX9074,WX9076,WX9078,WX9080,WX9082,
    WX9084,WX9536,WX9535,WX9538,WX9537,WX9540,WX9539,WX9542,WX9541,WX9544,
    WX9543,WX9546,WX9545,WX9548,WX9547,WX9550,WX9549,WX9552,WX9551,WX9554,
    WX9553,WX9556,WX9555,WX9558,WX9557,WX9560,WX9559,WX9562,WX9561,WX9564,
    WX9563,WX9566,WX9565,WX9568,WX9567,WX9570,WX9569,WX9572,WX9571,WX9574,
    WX9573,WX9576,WX9575,WX9578,WX9577,WX9580,WX9579,WX9582,WX9581,WX9584,
    WX9583,WX9586,WX9585,WX9588,WX9587,WX9590,WX9589,WX9592,WX9591,WX9594,
    WX9593,WX9596,WX9595,WX9598,WX9597,WX9696,WX9695,WX9698,WX9697,WX9700,
    WX9699,WX9702,WX9701,WX9704,WX9703,WX9706,WX9705,WX9708,WX9707,WX9710,
    WX9709,WX9712,WX9711,WX9714,WX9713,WX9716,WX9715,WX9718,WX9717,WX9720,
    WX9719,WX9722,WX9721,WX9724,WX9723,WX9726,WX9725,WX9728,WX9727,WX9730,
    WX9729,WX9732,WX9731,WX9734,WX9733,WX9736,WX9735,WX9738,WX9737,WX9740,
    WX9739,WX9742,WX9741,WX9744,WX9743,WX9746,WX9745,WX9748,WX9747,WX9750,
    WX9749,WX9752,WX9751,WX9754,WX9753,WX9756,WX9755,WX9758,WX9757,WX9760,
    WX9759,WX9762,WX9761,WX9764,WX9763,WX9766,WX9765,WX9768,WX9767,WX9770,
    WX9769,WX9772,WX9771,WX9774,WX9773,WX9776,WX9775,WX9778,WX9777,WX9780,
    WX9779,WX9782,WX9781,WX9784,WX9783,WX9786,WX9785,WX9788,WX9787,WX9790,
    WX9789,WX9792,WX9791,WX9794,WX9793,WX9796,WX9795,WX9798,WX9797,WX9800,
    WX9799,WX9802,WX9801,WX9804,WX9803,WX9806,WX9805,WX9808,WX9807,WX9810,
    WX9809,WX9812,WX9811,WX9814,WX9813,WX9816,WX9815,WX9818,WX9817,WX9820,
    WX9819,WX9822,WX9821,WX9824,WX9823,WX9826,WX9825,WX9828,WX9827,WX9830,
    WX9829,WX9832,WX9831,WX9834,WX9833,WX9836,WX9835,WX9838,WX9837,WX9840,
    WX9839,WX9842,WX9841,WX9844,WX9843,WX9846,WX9845,WX9848,WX9847,WX9850,
    WX9849,WX9852,WX9851,WX9854,WX9853,WX9856,WX9855,WX9858,WX9857,WX9860,
    WX9859,WX9862,WX9861,WX9864,WX9863,WX9866,WX9865,WX9868,WX9867,WX9870,
    WX9869,WX9872,WX9871,WX9874,WX9873,WX9876,WX9875,WX9878,WX9877,WX9880,
    WX9879,WX9882,WX9881,WX9884,WX9883,WX9886,WX9885,WX9888,WX9887,WX9890,
    WX9889,WX9892,WX9891,WX9894,WX9893,WX9896,WX9895,WX9898,WX9897,WX9900,
    WX9899,WX9902,WX9901,WX9904,WX9903,WX9906,WX9905,WX9908,WX9907,WX9910,
    WX9909,WX9912,WX9911,WX9914,WX9913,WX9916,WX9915,WX9918,WX9917,WX9920,
    WX9919,WX9922,WX9921,WX9924,WX9923,WX9926,WX9925,WX9928,WX9927,WX9930,
    WX9929,WX9932,WX9931,WX9934,WX9933,WX9936,WX9935,WX9938,WX9937,WX9940,
    WX9939,WX9942,WX9941,WX9944,WX9943,WX9946,WX9945,WX9948,WX9947,WX9950,
    WX9949,WX10315,WX10317,WX10319,WX10321,WX10323,WX10325,WX10327,WX10329,
    WX10331,WX10333,WX10335,WX10337,WX10339,WX10341,WX10343,WX10345,WX10347,
    WX10349,WX10351,WX10353,WX10355,WX10357,WX10359,WX10361,WX10363,WX10365,
    WX10367,WX10369,WX10371,WX10373,WX10375,WX10377,WX10829,WX10828,WX10831,
    WX10830,WX10833,WX10832,WX10835,WX10834,WX10837,WX10836,WX10839,WX10838,
    WX10841,WX10840,WX10843,WX10842,WX10845,WX10844,WX10847,WX10846,WX10849,
    WX10848,WX10851,WX10850,WX10853,WX10852,WX10855,WX10854,WX10857,WX10856,
    WX10859,WX10858,WX10861,WX10860,WX10863,WX10862,WX10865,WX10864,WX10867,
    WX10866,WX10869,WX10868,WX10871,WX10870,WX10873,WX10872,WX10875,WX10874,
    WX10877,WX10876,WX10879,WX10878,WX10881,WX10880,WX10883,WX10882,WX10885,
    WX10884,WX10887,WX10886,WX10889,WX10888,WX10891,WX10890,WX10989,WX10988,
    WX10991,WX10990,WX10993,WX10992,WX10995,WX10994,WX10997,WX10996,WX10999,
    WX10998,WX11001,WX11000,WX11003,WX11002,WX11005,WX11004,WX11007,WX11006,
    WX11009,WX11008,WX11011,WX11010,WX11013,WX11012,WX11015,WX11014,WX11017,
    WX11016,WX11019,WX11018,WX11021,WX11020,WX11023,WX11022,WX11025,WX11024,
    WX11027,WX11026,WX11029,WX11028,WX11031,WX11030,WX11033,WX11032,WX11035,
    WX11034,WX11037,WX11036,WX11039,WX11038,WX11041,WX11040,WX11043,WX11042,
    WX11045,WX11044,WX11047,WX11046,WX11049,WX11048,WX11051,WX11050,WX11053,
    WX11052,WX11055,WX11054,WX11057,WX11056,WX11059,WX11058,WX11061,WX11060,
    WX11063,WX11062,WX11065,WX11064,WX11067,WX11066,WX11069,WX11068,WX11071,
    WX11070,WX11073,WX11072,WX11075,WX11074,WX11077,WX11076,WX11079,WX11078,
    WX11081,WX11080,WX11083,WX11082,WX11085,WX11084,WX11087,WX11086,WX11089,
    WX11088,WX11091,WX11090,WX11093,WX11092,WX11095,WX11094,WX11097,WX11096,
    WX11099,WX11098,WX11101,WX11100,WX11103,WX11102,WX11105,WX11104,WX11107,
    WX11106,WX11109,WX11108,WX11111,WX11110,WX11113,WX11112,WX11115,WX11114,
    WX11117,WX11116,WX11119,WX11118,WX11121,WX11120,WX11123,WX11122,WX11125,
    WX11124,WX11127,WX11126,WX11129,WX11128,WX11131,WX11130,WX11133,WX11132,
    WX11135,WX11134,WX11137,WX11136,WX11139,WX11138,WX11141,WX11140,WX11143,
    WX11142,WX11145,WX11144,WX11147,WX11146,WX11149,WX11148,WX11151,WX11150,
    WX11153,WX11152,WX11155,WX11154,WX11157,WX11156,WX11159,WX11158,WX11161,
    WX11160,WX11163,WX11162,WX11165,WX11164,WX11167,WX11166,WX11169,WX11168,
    WX11171,WX11170,WX11173,WX11172,WX11175,WX11174,WX11177,WX11176,WX11179,
    WX11178,WX11181,WX11180,WX11183,WX11182,WX11185,WX11184,WX11187,WX11186,
    WX11189,WX11188,WX11191,WX11190,WX11193,WX11192,WX11195,WX11194,WX11197,
    WX11196,WX11199,WX11198,WX11201,WX11200,WX11203,WX11202,WX11205,WX11204,
    WX11207,WX11206,WX11209,WX11208,WX11211,WX11210,WX11213,WX11212,WX11215,
    WX11214,WX11217,WX11216,WX11219,WX11218,WX11221,WX11220,WX11223,WX11222,
    WX11225,WX11224,WX11227,WX11226,WX11229,WX11228,WX11231,WX11230,WX11233,
    WX11232,WX11235,WX11234,WX11237,WX11236,WX11239,WX11238,WX11241,WX11240,
    WX11243,WX11242,WX11608,WX11610,WX11612,WX11614,WX11616,WX11618,WX11620,
    WX11622,WX11624,WX11626,WX11628,WX11630,WX11632,WX11634,WX11636,WX11638,
    WX11640,WX11642,WX11644,WX11646,WX11648,WX11650,WX11652,WX11654,WX11656,
    WX11658,WX11660,WX11662,WX11664,WX11666,WX11668,WX11670,WX37,WX1003,WX41,
    WX1004,WX45,WX47,WX38,WX48,WX51,WX55,WX59,WX61,WX52,WX62,WX65,WX69,WX73,
    WX75,WX66,WX76,WX79,WX83,WX87,WX89,WX80,WX90,WX93,WX97,WX101,WX103,WX94,
    WX104,WX107,WX111,WX115,WX117,WX108,WX118,WX121,WX125,WX129,WX131,WX122,
    WX132,WX135,WX139,WX143,WX145,WX136,WX146,WX149,WX153,WX157,WX159,WX150,
    WX160,WX163,WX167,WX171,WX173,WX164,WX174,WX177,WX181,WX185,WX187,WX178,
    WX188,WX191,WX195,WX199,WX201,WX192,WX202,WX205,WX209,WX213,WX215,WX206,
    WX216,WX219,WX223,WX227,WX229,WX220,WX230,WX233,WX237,WX241,WX243,WX234,
    WX244,WX247,WX251,WX255,WX257,WX248,WX258,WX261,WX265,WX269,WX271,WX262,
    WX272,WX275,WX279,WX283,WX285,WX276,WX286,WX289,WX293,WX297,WX299,WX290,
    WX300,WX303,WX307,WX311,WX313,WX304,WX314,WX317,WX321,WX325,WX327,WX318,
    WX328,WX331,WX335,WX339,WX341,WX332,WX342,WX345,WX349,WX353,WX355,WX346,
    WX356,WX359,WX363,WX367,WX369,WX360,WX370,WX373,WX377,WX381,WX383,WX374,
    WX384,WX387,WX391,WX395,WX397,WX388,WX398,WX401,WX405,WX409,WX411,WX402,
    WX412,WX415,WX419,WX423,WX425,WX416,WX426,WX429,WX433,WX437,WX439,WX430,
    WX440,WX443,WX447,WX451,WX453,WX444,WX454,WX457,WX461,WX465,WX467,WX458,
    WX468,WX471,WX475,WX479,WX481,WX472,WX482,WX483,WX548,WX965,WX549,WX967,
    WX550,WX969,WX551,WX971,WX552,WX973,WX553,WX975,WX554,WX977,WX555,WX979,
    WX556,WX981,WX557,WX983,WX558,WX985,WX559,WX987,WX560,WX989,WX561,WX991,
    WX562,WX993,WX563,WX995,WX564,WX933,WX565,WX935,WX566,WX937,WX567,WX939,
    WX568,WX941,WX569,WX943,WX570,WX945,WX571,WX947,WX572,WX949,WX573,WX951,
    WX574,WX953,WX575,WX955,WX576,WX957,WX577,WX959,WX578,WX961,WX579,WX963,
    WX580,WX581,WX582,WX583,WX584,WX585,WX586,WX587,WX588,WX589,WX590,WX591,
    WX592,WX593,WX594,WX595,WX596,WX597,WX598,WX599,WX600,WX601,WX602,WX603,
    WX604,WX605,WX606,WX607,WX608,WX609,WX610,WX611,WX612,WX613,WX614,WX615,
    WX616,WX617,WX618,WX619,WX620,WX621,WX622,WX623,WX624,WX625,WX626,WX627,
    WX628,WX629,WX630,WX631,WX632,WX633,WX634,WX635,WX636,WX637,WX638,WX639,
    WX640,WX641,WX642,WX643,WX932,WX916,WX934,WX917,WX936,WX918,WX938,WX919,
    WX940,WX920,WX942,WX921,WX944,WX922,WX946,WX923,WX948,WX924,WX950,WX925,
    WX952,WX926,WX954,WX927,WX956,WX928,WX958,WX929,WX960,WX930,WX962,WX931,
    WX964,WX900,WX966,WX901,WX968,WX902,WX970,WX903,WX972,WX904,WX974,WX905,
    WX976,WX906,WX978,WX907,WX980,WX908,WX982,WX909,WX984,WX910,WX986,WX911,
    WX988,WX912,WX990,WX913,WX992,WX914,WX994,WX915,WX996,WX997,WX998,WX999,
    WX1000,WX1001,WX1002,WX1005,WX1009,WX1011,WX1010,WX1016,WX1018,WX1017,
    WX1023,WX1025,WX1024,WX1030,WX1032,WX1031,WX1037,WX1039,WX1038,WX1044,
    WX1046,WX1045,WX1051,WX1053,WX1052,WX1058,WX1060,WX1059,WX1065,WX1067,
    WX1066,WX1072,WX1074,WX1073,WX1079,WX1081,WX1080,WX1086,WX1088,WX1087,
    WX1093,WX1095,WX1094,WX1100,WX1102,WX1101,WX1107,WX1109,WX1108,WX1114,
    WX1116,WX1115,WX1121,WX1123,WX1122,WX1128,WX1130,WX1129,WX1135,WX1137,
    WX1136,WX1142,WX1144,WX1143,WX1149,WX1151,WX1150,WX1156,WX1158,WX1157,
    WX1163,WX1165,WX1164,WX1170,WX1172,WX1171,WX1177,WX1179,WX1178,WX1184,
    WX1186,WX1185,WX1191,WX1193,WX1192,WX1198,WX1200,WX1199,WX1205,WX1207,
    WX1206,WX1212,WX1214,WX1213,WX1219,WX1221,WX1220,WX1226,WX1228,WX1227,
    WX1230,WX1263,WX1330,WX2296,WX1334,WX2297,WX1338,WX1340,WX1331,WX1341,
    WX1344,WX1348,WX1352,WX1354,WX1345,WX1355,WX1358,WX1362,WX1366,WX1368,
    WX1359,WX1369,WX1372,WX1376,WX1380,WX1382,WX1373,WX1383,WX1386,WX1390,
    WX1394,WX1396,WX1387,WX1397,WX1400,WX1404,WX1408,WX1410,WX1401,WX1411,
    WX1414,WX1418,WX1422,WX1424,WX1415,WX1425,WX1428,WX1432,WX1436,WX1438,
    WX1429,WX1439,WX1442,WX1446,WX1450,WX1452,WX1443,WX1453,WX1456,WX1460,
    WX1464,WX1466,WX1457,WX1467,WX1470,WX1474,WX1478,WX1480,WX1471,WX1481,
    WX1484,WX1488,WX1492,WX1494,WX1485,WX1495,WX1498,WX1502,WX1506,WX1508,
    WX1499,WX1509,WX1512,WX1516,WX1520,WX1522,WX1513,WX1523,WX1526,WX1530,
    WX1534,WX1536,WX1527,WX1537,WX1540,WX1544,WX1548,WX1550,WX1541,WX1551,
    WX1554,WX1558,WX1562,WX1564,WX1555,WX1565,WX1568,WX1572,WX1576,WX1578,
    WX1569,WX1579,WX1582,WX1586,WX1590,WX1592,WX1583,WX1593,WX1596,WX1600,
    WX1604,WX1606,WX1597,WX1607,WX1610,WX1614,WX1618,WX1620,WX1611,WX1621,
    WX1624,WX1628,WX1632,WX1634,WX1625,WX1635,WX1638,WX1642,WX1646,WX1648,
    WX1639,WX1649,WX1652,WX1656,WX1660,WX1662,WX1653,WX1663,WX1666,WX1670,
    WX1674,WX1676,WX1667,WX1677,WX1680,WX1684,WX1688,WX1690,WX1681,WX1691,
    WX1694,WX1698,WX1702,WX1704,WX1695,WX1705,WX1708,WX1712,WX1716,WX1718,
    WX1709,WX1719,WX1722,WX1726,WX1730,WX1732,WX1723,WX1733,WX1736,WX1740,
    WX1744,WX1746,WX1737,WX1747,WX1750,WX1754,WX1758,WX1760,WX1751,WX1761,
    WX1764,WX1768,WX1772,WX1774,WX1765,WX1775,WX1776,WX1841,WX2258,WX1842,
    WX2260,WX1843,WX2262,WX1844,WX2264,WX1845,WX2266,WX1846,WX2268,WX1847,
    WX2270,WX1848,WX2272,WX1849,WX2274,WX1850,WX2276,WX1851,WX2278,WX1852,
    WX2280,WX1853,WX2282,WX1854,WX2284,WX1855,WX2286,WX1856,WX2288,WX1857,
    WX2226,WX1858,WX2228,WX1859,WX2230,WX1860,WX2232,WX1861,WX2234,WX1862,
    WX2236,WX1863,WX2238,WX1864,WX2240,WX1865,WX2242,WX1866,WX2244,WX1867,
    WX2246,WX1868,WX2248,WX1869,WX2250,WX1870,WX2252,WX1871,WX2254,WX1872,
    WX2256,WX1873,WX1874,WX1875,WX1876,WX1877,WX1878,WX1879,WX1880,WX1881,
    WX1882,WX1883,WX1884,WX1885,WX1886,WX1887,WX1888,WX1889,WX1890,WX1891,
    WX1892,WX1893,WX1894,WX1895,WX1896,WX1897,WX1898,WX1899,WX1900,WX1901,
    WX1902,WX1903,WX1904,WX1905,WX1906,WX1907,WX1908,WX1909,WX1910,WX1911,
    WX1912,WX1913,WX1914,WX1915,WX1916,WX1917,WX1918,WX1919,WX1920,WX1921,
    WX1922,WX1923,WX1924,WX1925,WX1926,WX1927,WX1928,WX1929,WX1930,WX1931,
    WX1932,WX1933,WX1934,WX1935,WX1936,WX2225,WX2209,WX2227,WX2210,WX2229,
    WX2211,WX2231,WX2212,WX2233,WX2213,WX2235,WX2214,WX2237,WX2215,WX2239,
    WX2216,WX2241,WX2217,WX2243,WX2218,WX2245,WX2219,WX2247,WX2220,WX2249,
    WX2221,WX2251,WX2222,WX2253,WX2223,WX2255,WX2224,WX2257,WX2193,WX2259,
    WX2194,WX2261,WX2195,WX2263,WX2196,WX2265,WX2197,WX2267,WX2198,WX2269,
    WX2199,WX2271,WX2200,WX2273,WX2201,WX2275,WX2202,WX2277,WX2203,WX2279,
    WX2204,WX2281,WX2205,WX2283,WX2206,WX2285,WX2207,WX2287,WX2208,WX2289,
    WX2290,WX2291,WX2292,WX2293,WX2294,WX2295,WX2298,WX2302,WX2304,WX2303,
    WX2305,WX2309,WX2311,WX2310,WX2312,WX2316,WX2318,WX2317,WX2319,WX2323,
    WX2325,WX2324,WX2326,WX2330,WX2332,WX2331,WX2333,WX2337,WX2339,WX2338,
    WX2340,WX2344,WX2346,WX2345,WX2347,WX2351,WX2353,WX2352,WX2354,WX2358,
    WX2360,WX2359,WX2361,WX2365,WX2367,WX2366,WX2368,WX2372,WX2374,WX2373,
    WX2375,WX2379,WX2381,WX2380,WX2382,WX2386,WX2388,WX2387,WX2389,WX2393,
    WX2395,WX2394,WX2396,WX2400,WX2402,WX2401,WX2403,WX2407,WX2409,WX2408,
    WX2410,WX2414,WX2416,WX2415,WX2417,WX2421,WX2423,WX2422,WX2424,WX2428,
    WX2430,WX2429,WX2431,WX2435,WX2437,WX2436,WX2438,WX2442,WX2444,WX2443,
    WX2445,WX2449,WX2451,WX2450,WX2452,WX2456,WX2458,WX2457,WX2459,WX2463,
    WX2465,WX2464,WX2466,WX2470,WX2472,WX2471,WX2473,WX2477,WX2479,WX2478,
    WX2480,WX2484,WX2486,WX2485,WX2487,WX2491,WX2493,WX2492,WX2494,WX2498,
    WX2500,WX2499,WX2501,WX2505,WX2507,WX2506,WX2508,WX2512,WX2514,WX2513,
    WX2515,WX2519,WX2521,WX2520,WX2522,WX2523,WX2556,WX2623,WX3589,WX2627,
    WX3590,WX2631,WX2633,WX2624,WX2634,WX2637,WX2641,WX2645,WX2647,WX2638,
    WX2648,WX2651,WX2655,WX2659,WX2661,WX2652,WX2662,WX2665,WX2669,WX2673,
    WX2675,WX2666,WX2676,WX2679,WX2683,WX2687,WX2689,WX2680,WX2690,WX2693,
    WX2697,WX2701,WX2703,WX2694,WX2704,WX2707,WX2711,WX2715,WX2717,WX2708,
    WX2718,WX2721,WX2725,WX2729,WX2731,WX2722,WX2732,WX2735,WX2739,WX2743,
    WX2745,WX2736,WX2746,WX2749,WX2753,WX2757,WX2759,WX2750,WX2760,WX2763,
    WX2767,WX2771,WX2773,WX2764,WX2774,WX2777,WX2781,WX2785,WX2787,WX2778,
    WX2788,WX2791,WX2795,WX2799,WX2801,WX2792,WX2802,WX2805,WX2809,WX2813,
    WX2815,WX2806,WX2816,WX2819,WX2823,WX2827,WX2829,WX2820,WX2830,WX2833,
    WX2837,WX2841,WX2843,WX2834,WX2844,WX2847,WX2851,WX2855,WX2857,WX2848,
    WX2858,WX2861,WX2865,WX2869,WX2871,WX2862,WX2872,WX2875,WX2879,WX2883,
    WX2885,WX2876,WX2886,WX2889,WX2893,WX2897,WX2899,WX2890,WX2900,WX2903,
    WX2907,WX2911,WX2913,WX2904,WX2914,WX2917,WX2921,WX2925,WX2927,WX2918,
    WX2928,WX2931,WX2935,WX2939,WX2941,WX2932,WX2942,WX2945,WX2949,WX2953,
    WX2955,WX2946,WX2956,WX2959,WX2963,WX2967,WX2969,WX2960,WX2970,WX2973,
    WX2977,WX2981,WX2983,WX2974,WX2984,WX2987,WX2991,WX2995,WX2997,WX2988,
    WX2998,WX3001,WX3005,WX3009,WX3011,WX3002,WX3012,WX3015,WX3019,WX3023,
    WX3025,WX3016,WX3026,WX3029,WX3033,WX3037,WX3039,WX3030,WX3040,WX3043,
    WX3047,WX3051,WX3053,WX3044,WX3054,WX3057,WX3061,WX3065,WX3067,WX3058,
    WX3068,WX3069,WX3134,WX3551,WX3135,WX3553,WX3136,WX3555,WX3137,WX3557,
    WX3138,WX3559,WX3139,WX3561,WX3140,WX3563,WX3141,WX3565,WX3142,WX3567,
    WX3143,WX3569,WX3144,WX3571,WX3145,WX3573,WX3146,WX3575,WX3147,WX3577,
    WX3148,WX3579,WX3149,WX3581,WX3150,WX3519,WX3151,WX3521,WX3152,WX3523,
    WX3153,WX3525,WX3154,WX3527,WX3155,WX3529,WX3156,WX3531,WX3157,WX3533,
    WX3158,WX3535,WX3159,WX3537,WX3160,WX3539,WX3161,WX3541,WX3162,WX3543,
    WX3163,WX3545,WX3164,WX3547,WX3165,WX3549,WX3166,WX3167,WX3168,WX3169,
    WX3170,WX3171,WX3172,WX3173,WX3174,WX3175,WX3176,WX3177,WX3178,WX3179,
    WX3180,WX3181,WX3182,WX3183,WX3184,WX3185,WX3186,WX3187,WX3188,WX3189,
    WX3190,WX3191,WX3192,WX3193,WX3194,WX3195,WX3196,WX3197,WX3198,WX3199,
    WX3200,WX3201,WX3202,WX3203,WX3204,WX3205,WX3206,WX3207,WX3208,WX3209,
    WX3210,WX3211,WX3212,WX3213,WX3214,WX3215,WX3216,WX3217,WX3218,WX3219,
    WX3220,WX3221,WX3222,WX3223,WX3224,WX3225,WX3226,WX3227,WX3228,WX3229,
    WX3518,WX3502,WX3520,WX3503,WX3522,WX3504,WX3524,WX3505,WX3526,WX3506,
    WX3528,WX3507,WX3530,WX3508,WX3532,WX3509,WX3534,WX3510,WX3536,WX3511,
    WX3538,WX3512,WX3540,WX3513,WX3542,WX3514,WX3544,WX3515,WX3546,WX3516,
    WX3548,WX3517,WX3550,WX3486,WX3552,WX3487,WX3554,WX3488,WX3556,WX3489,
    WX3558,WX3490,WX3560,WX3491,WX3562,WX3492,WX3564,WX3493,WX3566,WX3494,
    WX3568,WX3495,WX3570,WX3496,WX3572,WX3497,WX3574,WX3498,WX3576,WX3499,
    WX3578,WX3500,WX3580,WX3501,WX3582,WX3583,WX3584,WX3585,WX3586,WX3587,
    WX3588,WX3591,WX3595,WX3597,WX3596,WX3598,WX3602,WX3604,WX3603,WX3605,
    WX3609,WX3611,WX3610,WX3612,WX3616,WX3618,WX3617,WX3619,WX3623,WX3625,
    WX3624,WX3626,WX3630,WX3632,WX3631,WX3633,WX3637,WX3639,WX3638,WX3640,
    WX3644,WX3646,WX3645,WX3647,WX3651,WX3653,WX3652,WX3654,WX3658,WX3660,
    WX3659,WX3661,WX3665,WX3667,WX3666,WX3668,WX3672,WX3674,WX3673,WX3675,
    WX3679,WX3681,WX3680,WX3682,WX3686,WX3688,WX3687,WX3689,WX3693,WX3695,
    WX3694,WX3696,WX3700,WX3702,WX3701,WX3703,WX3707,WX3709,WX3708,WX3710,
    WX3714,WX3716,WX3715,WX3717,WX3721,WX3723,WX3722,WX3724,WX3728,WX3730,
    WX3729,WX3731,WX3735,WX3737,WX3736,WX3738,WX3742,WX3744,WX3743,WX3745,
    WX3749,WX3751,WX3750,WX3752,WX3756,WX3758,WX3757,WX3759,WX3763,WX3765,
    WX3764,WX3766,WX3770,WX3772,WX3771,WX3773,WX3777,WX3779,WX3778,WX3780,
    WX3784,WX3786,WX3785,WX3787,WX3791,WX3793,WX3792,WX3794,WX3798,WX3800,
    WX3799,WX3801,WX3805,WX3807,WX3806,WX3808,WX3812,WX3814,WX3813,WX3815,
    WX3816,WX3849,WX3916,WX4882,WX3920,WX4883,WX3924,WX3926,WX3917,WX3927,
    WX3930,WX3934,WX3938,WX3940,WX3931,WX3941,WX3944,WX3948,WX3952,WX3954,
    WX3945,WX3955,WX3958,WX3962,WX3966,WX3968,WX3959,WX3969,WX3972,WX3976,
    WX3980,WX3982,WX3973,WX3983,WX3986,WX3990,WX3994,WX3996,WX3987,WX3997,
    WX4000,WX4004,WX4008,WX4010,WX4001,WX4011,WX4014,WX4018,WX4022,WX4024,
    WX4015,WX4025,WX4028,WX4032,WX4036,WX4038,WX4029,WX4039,WX4042,WX4046,
    WX4050,WX4052,WX4043,WX4053,WX4056,WX4060,WX4064,WX4066,WX4057,WX4067,
    WX4070,WX4074,WX4078,WX4080,WX4071,WX4081,WX4084,WX4088,WX4092,WX4094,
    WX4085,WX4095,WX4098,WX4102,WX4106,WX4108,WX4099,WX4109,WX4112,WX4116,
    WX4120,WX4122,WX4113,WX4123,WX4126,WX4130,WX4134,WX4136,WX4127,WX4137,
    WX4140,WX4144,WX4148,WX4150,WX4141,WX4151,WX4154,WX4158,WX4162,WX4164,
    WX4155,WX4165,WX4168,WX4172,WX4176,WX4178,WX4169,WX4179,WX4182,WX4186,
    WX4190,WX4192,WX4183,WX4193,WX4196,WX4200,WX4204,WX4206,WX4197,WX4207,
    WX4210,WX4214,WX4218,WX4220,WX4211,WX4221,WX4224,WX4228,WX4232,WX4234,
    WX4225,WX4235,WX4238,WX4242,WX4246,WX4248,WX4239,WX4249,WX4252,WX4256,
    WX4260,WX4262,WX4253,WX4263,WX4266,WX4270,WX4274,WX4276,WX4267,WX4277,
    WX4280,WX4284,WX4288,WX4290,WX4281,WX4291,WX4294,WX4298,WX4302,WX4304,
    WX4295,WX4305,WX4308,WX4312,WX4316,WX4318,WX4309,WX4319,WX4322,WX4326,
    WX4330,WX4332,WX4323,WX4333,WX4336,WX4340,WX4344,WX4346,WX4337,WX4347,
    WX4350,WX4354,WX4358,WX4360,WX4351,WX4361,WX4362,WX4427,WX4844,WX4428,
    WX4846,WX4429,WX4848,WX4430,WX4850,WX4431,WX4852,WX4432,WX4854,WX4433,
    WX4856,WX4434,WX4858,WX4435,WX4860,WX4436,WX4862,WX4437,WX4864,WX4438,
    WX4866,WX4439,WX4868,WX4440,WX4870,WX4441,WX4872,WX4442,WX4874,WX4443,
    WX4812,WX4444,WX4814,WX4445,WX4816,WX4446,WX4818,WX4447,WX4820,WX4448,
    WX4822,WX4449,WX4824,WX4450,WX4826,WX4451,WX4828,WX4452,WX4830,WX4453,
    WX4832,WX4454,WX4834,WX4455,WX4836,WX4456,WX4838,WX4457,WX4840,WX4458,
    WX4842,WX4459,WX4460,WX4461,WX4462,WX4463,WX4464,WX4465,WX4466,WX4467,
    WX4468,WX4469,WX4470,WX4471,WX4472,WX4473,WX4474,WX4475,WX4476,WX4477,
    WX4478,WX4479,WX4480,WX4481,WX4482,WX4483,WX4484,WX4485,WX4486,WX4487,
    WX4488,WX4489,WX4490,WX4491,WX4492,WX4493,WX4494,WX4495,WX4496,WX4497,
    WX4498,WX4499,WX4500,WX4501,WX4502,WX4503,WX4504,WX4505,WX4506,WX4507,
    WX4508,WX4509,WX4510,WX4511,WX4512,WX4513,WX4514,WX4515,WX4516,WX4517,
    WX4518,WX4519,WX4520,WX4521,WX4522,WX4811,WX4795,WX4813,WX4796,WX4815,
    WX4797,WX4817,WX4798,WX4819,WX4799,WX4821,WX4800,WX4823,WX4801,WX4825,
    WX4802,WX4827,WX4803,WX4829,WX4804,WX4831,WX4805,WX4833,WX4806,WX4835,
    WX4807,WX4837,WX4808,WX4839,WX4809,WX4841,WX4810,WX4843,WX4779,WX4845,
    WX4780,WX4847,WX4781,WX4849,WX4782,WX4851,WX4783,WX4853,WX4784,WX4855,
    WX4785,WX4857,WX4786,WX4859,WX4787,WX4861,WX4788,WX4863,WX4789,WX4865,
    WX4790,WX4867,WX4791,WX4869,WX4792,WX4871,WX4793,WX4873,WX4794,WX4875,
    WX4876,WX4877,WX4878,WX4879,WX4880,WX4881,WX4884,WX4888,WX4890,WX4889,
    WX4891,WX4895,WX4897,WX4896,WX4898,WX4902,WX4904,WX4903,WX4905,WX4909,
    WX4911,WX4910,WX4912,WX4916,WX4918,WX4917,WX4919,WX4923,WX4925,WX4924,
    WX4926,WX4930,WX4932,WX4931,WX4933,WX4937,WX4939,WX4938,WX4940,WX4944,
    WX4946,WX4945,WX4947,WX4951,WX4953,WX4952,WX4954,WX4958,WX4960,WX4959,
    WX4961,WX4965,WX4967,WX4966,WX4968,WX4972,WX4974,WX4973,WX4975,WX4979,
    WX4981,WX4980,WX4982,WX4986,WX4988,WX4987,WX4989,WX4993,WX4995,WX4994,
    WX4996,WX5000,WX5002,WX5001,WX5003,WX5007,WX5009,WX5008,WX5010,WX5014,
    WX5016,WX5015,WX5017,WX5021,WX5023,WX5022,WX5024,WX5028,WX5030,WX5029,
    WX5031,WX5035,WX5037,WX5036,WX5038,WX5042,WX5044,WX5043,WX5045,WX5049,
    WX5051,WX5050,WX5052,WX5056,WX5058,WX5057,WX5059,WX5063,WX5065,WX5064,
    WX5066,WX5070,WX5072,WX5071,WX5073,WX5077,WX5079,WX5078,WX5080,WX5084,
    WX5086,WX5085,WX5087,WX5091,WX5093,WX5092,WX5094,WX5098,WX5100,WX5099,
    WX5101,WX5105,WX5107,WX5106,WX5108,WX5109,WX5142,WX5209,WX6175,WX5213,
    WX6176,WX5217,WX5219,WX5210,WX5220,WX5223,WX5227,WX5231,WX5233,WX5224,
    WX5234,WX5237,WX5241,WX5245,WX5247,WX5238,WX5248,WX5251,WX5255,WX5259,
    WX5261,WX5252,WX5262,WX5265,WX5269,WX5273,WX5275,WX5266,WX5276,WX5279,
    WX5283,WX5287,WX5289,WX5280,WX5290,WX5293,WX5297,WX5301,WX5303,WX5294,
    WX5304,WX5307,WX5311,WX5315,WX5317,WX5308,WX5318,WX5321,WX5325,WX5329,
    WX5331,WX5322,WX5332,WX5335,WX5339,WX5343,WX5345,WX5336,WX5346,WX5349,
    WX5353,WX5357,WX5359,WX5350,WX5360,WX5363,WX5367,WX5371,WX5373,WX5364,
    WX5374,WX5377,WX5381,WX5385,WX5387,WX5378,WX5388,WX5391,WX5395,WX5399,
    WX5401,WX5392,WX5402,WX5405,WX5409,WX5413,WX5415,WX5406,WX5416,WX5419,
    WX5423,WX5427,WX5429,WX5420,WX5430,WX5433,WX5437,WX5441,WX5443,WX5434,
    WX5444,WX5447,WX5451,WX5455,WX5457,WX5448,WX5458,WX5461,WX5465,WX5469,
    WX5471,WX5462,WX5472,WX5475,WX5479,WX5483,WX5485,WX5476,WX5486,WX5489,
    WX5493,WX5497,WX5499,WX5490,WX5500,WX5503,WX5507,WX5511,WX5513,WX5504,
    WX5514,WX5517,WX5521,WX5525,WX5527,WX5518,WX5528,WX5531,WX5535,WX5539,
    WX5541,WX5532,WX5542,WX5545,WX5549,WX5553,WX5555,WX5546,WX5556,WX5559,
    WX5563,WX5567,WX5569,WX5560,WX5570,WX5573,WX5577,WX5581,WX5583,WX5574,
    WX5584,WX5587,WX5591,WX5595,WX5597,WX5588,WX5598,WX5601,WX5605,WX5609,
    WX5611,WX5602,WX5612,WX5615,WX5619,WX5623,WX5625,WX5616,WX5626,WX5629,
    WX5633,WX5637,WX5639,WX5630,WX5640,WX5643,WX5647,WX5651,WX5653,WX5644,
    WX5654,WX5655,WX5720,WX6137,WX5721,WX6139,WX5722,WX6141,WX5723,WX6143,
    WX5724,WX6145,WX5725,WX6147,WX5726,WX6149,WX5727,WX6151,WX5728,WX6153,
    WX5729,WX6155,WX5730,WX6157,WX5731,WX6159,WX5732,WX6161,WX5733,WX6163,
    WX5734,WX6165,WX5735,WX6167,WX5736,WX6105,WX5737,WX6107,WX5738,WX6109,
    WX5739,WX6111,WX5740,WX6113,WX5741,WX6115,WX5742,WX6117,WX5743,WX6119,
    WX5744,WX6121,WX5745,WX6123,WX5746,WX6125,WX5747,WX6127,WX5748,WX6129,
    WX5749,WX6131,WX5750,WX6133,WX5751,WX6135,WX5752,WX5753,WX5754,WX5755,
    WX5756,WX5757,WX5758,WX5759,WX5760,WX5761,WX5762,WX5763,WX5764,WX5765,
    WX5766,WX5767,WX5768,WX5769,WX5770,WX5771,WX5772,WX5773,WX5774,WX5775,
    WX5776,WX5777,WX5778,WX5779,WX5780,WX5781,WX5782,WX5783,WX5784,WX5785,
    WX5786,WX5787,WX5788,WX5789,WX5790,WX5791,WX5792,WX5793,WX5794,WX5795,
    WX5796,WX5797,WX5798,WX5799,WX5800,WX5801,WX5802,WX5803,WX5804,WX5805,
    WX5806,WX5807,WX5808,WX5809,WX5810,WX5811,WX5812,WX5813,WX5814,WX5815,
    WX6104,WX6088,WX6106,WX6089,WX6108,WX6090,WX6110,WX6091,WX6112,WX6092,
    WX6114,WX6093,WX6116,WX6094,WX6118,WX6095,WX6120,WX6096,WX6122,WX6097,
    WX6124,WX6098,WX6126,WX6099,WX6128,WX6100,WX6130,WX6101,WX6132,WX6102,
    WX6134,WX6103,WX6136,WX6072,WX6138,WX6073,WX6140,WX6074,WX6142,WX6075,
    WX6144,WX6076,WX6146,WX6077,WX6148,WX6078,WX6150,WX6079,WX6152,WX6080,
    WX6154,WX6081,WX6156,WX6082,WX6158,WX6083,WX6160,WX6084,WX6162,WX6085,
    WX6164,WX6086,WX6166,WX6087,WX6168,WX6169,WX6170,WX6171,WX6172,WX6173,
    WX6174,WX6177,WX6181,WX6183,WX6182,WX6184,WX6188,WX6190,WX6189,WX6191,
    WX6195,WX6197,WX6196,WX6198,WX6202,WX6204,WX6203,WX6205,WX6209,WX6211,
    WX6210,WX6212,WX6216,WX6218,WX6217,WX6219,WX6223,WX6225,WX6224,WX6226,
    WX6230,WX6232,WX6231,WX6233,WX6237,WX6239,WX6238,WX6240,WX6244,WX6246,
    WX6245,WX6247,WX6251,WX6253,WX6252,WX6254,WX6258,WX6260,WX6259,WX6261,
    WX6265,WX6267,WX6266,WX6268,WX6272,WX6274,WX6273,WX6275,WX6279,WX6281,
    WX6280,WX6282,WX6286,WX6288,WX6287,WX6289,WX6293,WX6295,WX6294,WX6296,
    WX6300,WX6302,WX6301,WX6303,WX6307,WX6309,WX6308,WX6310,WX6314,WX6316,
    WX6315,WX6317,WX6321,WX6323,WX6322,WX6324,WX6328,WX6330,WX6329,WX6331,
    WX6335,WX6337,WX6336,WX6338,WX6342,WX6344,WX6343,WX6345,WX6349,WX6351,
    WX6350,WX6352,WX6356,WX6358,WX6357,WX6359,WX6363,WX6365,WX6364,WX6366,
    WX6370,WX6372,WX6371,WX6373,WX6377,WX6379,WX6378,WX6380,WX6384,WX6386,
    WX6385,WX6387,WX6391,WX6393,WX6392,WX6394,WX6398,WX6400,WX6399,WX6401,
    WX6402,WX6435,WX6502,WX7468,WX6506,WX7469,WX6510,WX6512,WX6503,WX6513,
    WX6516,WX6520,WX6524,WX6526,WX6517,WX6527,WX6530,WX6534,WX6538,WX6540,
    WX6531,WX6541,WX6544,WX6548,WX6552,WX6554,WX6545,WX6555,WX6558,WX6562,
    WX6566,WX6568,WX6559,WX6569,WX6572,WX6576,WX6580,WX6582,WX6573,WX6583,
    WX6586,WX6590,WX6594,WX6596,WX6587,WX6597,WX6600,WX6604,WX6608,WX6610,
    WX6601,WX6611,WX6614,WX6618,WX6622,WX6624,WX6615,WX6625,WX6628,WX6632,
    WX6636,WX6638,WX6629,WX6639,WX6642,WX6646,WX6650,WX6652,WX6643,WX6653,
    WX6656,WX6660,WX6664,WX6666,WX6657,WX6667,WX6670,WX6674,WX6678,WX6680,
    WX6671,WX6681,WX6684,WX6688,WX6692,WX6694,WX6685,WX6695,WX6698,WX6702,
    WX6706,WX6708,WX6699,WX6709,WX6712,WX6716,WX6720,WX6722,WX6713,WX6723,
    WX6726,WX6730,WX6734,WX6736,WX6727,WX6737,WX6740,WX6744,WX6748,WX6750,
    WX6741,WX6751,WX6754,WX6758,WX6762,WX6764,WX6755,WX6765,WX6768,WX6772,
    WX6776,WX6778,WX6769,WX6779,WX6782,WX6786,WX6790,WX6792,WX6783,WX6793,
    WX6796,WX6800,WX6804,WX6806,WX6797,WX6807,WX6810,WX6814,WX6818,WX6820,
    WX6811,WX6821,WX6824,WX6828,WX6832,WX6834,WX6825,WX6835,WX6838,WX6842,
    WX6846,WX6848,WX6839,WX6849,WX6852,WX6856,WX6860,WX6862,WX6853,WX6863,
    WX6866,WX6870,WX6874,WX6876,WX6867,WX6877,WX6880,WX6884,WX6888,WX6890,
    WX6881,WX6891,WX6894,WX6898,WX6902,WX6904,WX6895,WX6905,WX6908,WX6912,
    WX6916,WX6918,WX6909,WX6919,WX6922,WX6926,WX6930,WX6932,WX6923,WX6933,
    WX6936,WX6940,WX6944,WX6946,WX6937,WX6947,WX6948,WX7013,WX7430,WX7014,
    WX7432,WX7015,WX7434,WX7016,WX7436,WX7017,WX7438,WX7018,WX7440,WX7019,
    WX7442,WX7020,WX7444,WX7021,WX7446,WX7022,WX7448,WX7023,WX7450,WX7024,
    WX7452,WX7025,WX7454,WX7026,WX7456,WX7027,WX7458,WX7028,WX7460,WX7029,
    WX7398,WX7030,WX7400,WX7031,WX7402,WX7032,WX7404,WX7033,WX7406,WX7034,
    WX7408,WX7035,WX7410,WX7036,WX7412,WX7037,WX7414,WX7038,WX7416,WX7039,
    WX7418,WX7040,WX7420,WX7041,WX7422,WX7042,WX7424,WX7043,WX7426,WX7044,
    WX7428,WX7045,WX7046,WX7047,WX7048,WX7049,WX7050,WX7051,WX7052,WX7053,
    WX7054,WX7055,WX7056,WX7057,WX7058,WX7059,WX7060,WX7061,WX7062,WX7063,
    WX7064,WX7065,WX7066,WX7067,WX7068,WX7069,WX7070,WX7071,WX7072,WX7073,
    WX7074,WX7075,WX7076,WX7077,WX7078,WX7079,WX7080,WX7081,WX7082,WX7083,
    WX7084,WX7085,WX7086,WX7087,WX7088,WX7089,WX7090,WX7091,WX7092,WX7093,
    WX7094,WX7095,WX7096,WX7097,WX7098,WX7099,WX7100,WX7101,WX7102,WX7103,
    WX7104,WX7105,WX7106,WX7107,WX7108,WX7397,WX7381,WX7399,WX7382,WX7401,
    WX7383,WX7403,WX7384,WX7405,WX7385,WX7407,WX7386,WX7409,WX7387,WX7411,
    WX7388,WX7413,WX7389,WX7415,WX7390,WX7417,WX7391,WX7419,WX7392,WX7421,
    WX7393,WX7423,WX7394,WX7425,WX7395,WX7427,WX7396,WX7429,WX7365,WX7431,
    WX7366,WX7433,WX7367,WX7435,WX7368,WX7437,WX7369,WX7439,WX7370,WX7441,
    WX7371,WX7443,WX7372,WX7445,WX7373,WX7447,WX7374,WX7449,WX7375,WX7451,
    WX7376,WX7453,WX7377,WX7455,WX7378,WX7457,WX7379,WX7459,WX7380,WX7461,
    WX7462,WX7463,WX7464,WX7465,WX7466,WX7467,WX7470,WX7474,WX7476,WX7475,
    WX7477,WX7481,WX7483,WX7482,WX7484,WX7488,WX7490,WX7489,WX7491,WX7495,
    WX7497,WX7496,WX7498,WX7502,WX7504,WX7503,WX7505,WX7509,WX7511,WX7510,
    WX7512,WX7516,WX7518,WX7517,WX7519,WX7523,WX7525,WX7524,WX7526,WX7530,
    WX7532,WX7531,WX7533,WX7537,WX7539,WX7538,WX7540,WX7544,WX7546,WX7545,
    WX7547,WX7551,WX7553,WX7552,WX7554,WX7558,WX7560,WX7559,WX7561,WX7565,
    WX7567,WX7566,WX7568,WX7572,WX7574,WX7573,WX7575,WX7579,WX7581,WX7580,
    WX7582,WX7586,WX7588,WX7587,WX7589,WX7593,WX7595,WX7594,WX7596,WX7600,
    WX7602,WX7601,WX7603,WX7607,WX7609,WX7608,WX7610,WX7614,WX7616,WX7615,
    WX7617,WX7621,WX7623,WX7622,WX7624,WX7628,WX7630,WX7629,WX7631,WX7635,
    WX7637,WX7636,WX7638,WX7642,WX7644,WX7643,WX7645,WX7649,WX7651,WX7650,
    WX7652,WX7656,WX7658,WX7657,WX7659,WX7663,WX7665,WX7664,WX7666,WX7670,
    WX7672,WX7671,WX7673,WX7677,WX7679,WX7678,WX7680,WX7684,WX7686,WX7685,
    WX7687,WX7691,WX7693,WX7692,WX7694,WX7695,WX7728,WX7795,WX8761,WX7799,
    WX8762,WX7803,WX7805,WX7796,WX7806,WX7809,WX7813,WX7817,WX7819,WX7810,
    WX7820,WX7823,WX7827,WX7831,WX7833,WX7824,WX7834,WX7837,WX7841,WX7845,
    WX7847,WX7838,WX7848,WX7851,WX7855,WX7859,WX7861,WX7852,WX7862,WX7865,
    WX7869,WX7873,WX7875,WX7866,WX7876,WX7879,WX7883,WX7887,WX7889,WX7880,
    WX7890,WX7893,WX7897,WX7901,WX7903,WX7894,WX7904,WX7907,WX7911,WX7915,
    WX7917,WX7908,WX7918,WX7921,WX7925,WX7929,WX7931,WX7922,WX7932,WX7935,
    WX7939,WX7943,WX7945,WX7936,WX7946,WX7949,WX7953,WX7957,WX7959,WX7950,
    WX7960,WX7963,WX7967,WX7971,WX7973,WX7964,WX7974,WX7977,WX7981,WX7985,
    WX7987,WX7978,WX7988,WX7991,WX7995,WX7999,WX8001,WX7992,WX8002,WX8005,
    WX8009,WX8013,WX8015,WX8006,WX8016,WX8019,WX8023,WX8027,WX8029,WX8020,
    WX8030,WX8033,WX8037,WX8041,WX8043,WX8034,WX8044,WX8047,WX8051,WX8055,
    WX8057,WX8048,WX8058,WX8061,WX8065,WX8069,WX8071,WX8062,WX8072,WX8075,
    WX8079,WX8083,WX8085,WX8076,WX8086,WX8089,WX8093,WX8097,WX8099,WX8090,
    WX8100,WX8103,WX8107,WX8111,WX8113,WX8104,WX8114,WX8117,WX8121,WX8125,
    WX8127,WX8118,WX8128,WX8131,WX8135,WX8139,WX8141,WX8132,WX8142,WX8145,
    WX8149,WX8153,WX8155,WX8146,WX8156,WX8159,WX8163,WX8167,WX8169,WX8160,
    WX8170,WX8173,WX8177,WX8181,WX8183,WX8174,WX8184,WX8187,WX8191,WX8195,
    WX8197,WX8188,WX8198,WX8201,WX8205,WX8209,WX8211,WX8202,WX8212,WX8215,
    WX8219,WX8223,WX8225,WX8216,WX8226,WX8229,WX8233,WX8237,WX8239,WX8230,
    WX8240,WX8241,WX8306,WX8723,WX8307,WX8725,WX8308,WX8727,WX8309,WX8729,
    WX8310,WX8731,WX8311,WX8733,WX8312,WX8735,WX8313,WX8737,WX8314,WX8739,
    WX8315,WX8741,WX8316,WX8743,WX8317,WX8745,WX8318,WX8747,WX8319,WX8749,
    WX8320,WX8751,WX8321,WX8753,WX8322,WX8691,WX8323,WX8693,WX8324,WX8695,
    WX8325,WX8697,WX8326,WX8699,WX8327,WX8701,WX8328,WX8703,WX8329,WX8705,
    WX8330,WX8707,WX8331,WX8709,WX8332,WX8711,WX8333,WX8713,WX8334,WX8715,
    WX8335,WX8717,WX8336,WX8719,WX8337,WX8721,WX8338,WX8339,WX8340,WX8341,
    WX8342,WX8343,WX8344,WX8345,WX8346,WX8347,WX8348,WX8349,WX8350,WX8351,
    WX8352,WX8353,WX8354,WX8355,WX8356,WX8357,WX8358,WX8359,WX8360,WX8361,
    WX8362,WX8363,WX8364,WX8365,WX8366,WX8367,WX8368,WX8369,WX8370,WX8371,
    WX8372,WX8373,WX8374,WX8375,WX8376,WX8377,WX8378,WX8379,WX8380,WX8381,
    WX8382,WX8383,WX8384,WX8385,WX8386,WX8387,WX8388,WX8389,WX8390,WX8391,
    WX8392,WX8393,WX8394,WX8395,WX8396,WX8397,WX8398,WX8399,WX8400,WX8401,
    WX8690,WX8674,WX8692,WX8675,WX8694,WX8676,WX8696,WX8677,WX8698,WX8678,
    WX8700,WX8679,WX8702,WX8680,WX8704,WX8681,WX8706,WX8682,WX8708,WX8683,
    WX8710,WX8684,WX8712,WX8685,WX8714,WX8686,WX8716,WX8687,WX8718,WX8688,
    WX8720,WX8689,WX8722,WX8658,WX8724,WX8659,WX8726,WX8660,WX8728,WX8661,
    WX8730,WX8662,WX8732,WX8663,WX8734,WX8664,WX8736,WX8665,WX8738,WX8666,
    WX8740,WX8667,WX8742,WX8668,WX8744,WX8669,WX8746,WX8670,WX8748,WX8671,
    WX8750,WX8672,WX8752,WX8673,WX8754,WX8755,WX8756,WX8757,WX8758,WX8759,
    WX8760,WX8763,WX8767,WX8769,WX8768,WX8770,WX8774,WX8776,WX8775,WX8777,
    WX8781,WX8783,WX8782,WX8784,WX8788,WX8790,WX8789,WX8791,WX8795,WX8797,
    WX8796,WX8798,WX8802,WX8804,WX8803,WX8805,WX8809,WX8811,WX8810,WX8812,
    WX8816,WX8818,WX8817,WX8819,WX8823,WX8825,WX8824,WX8826,WX8830,WX8832,
    WX8831,WX8833,WX8837,WX8839,WX8838,WX8840,WX8844,WX8846,WX8845,WX8847,
    WX8851,WX8853,WX8852,WX8854,WX8858,WX8860,WX8859,WX8861,WX8865,WX8867,
    WX8866,WX8868,WX8872,WX8874,WX8873,WX8875,WX8879,WX8881,WX8880,WX8882,
    WX8886,WX8888,WX8887,WX8889,WX8893,WX8895,WX8894,WX8896,WX8900,WX8902,
    WX8901,WX8903,WX8907,WX8909,WX8908,WX8910,WX8914,WX8916,WX8915,WX8917,
    WX8921,WX8923,WX8922,WX8924,WX8928,WX8930,WX8929,WX8931,WX8935,WX8937,
    WX8936,WX8938,WX8942,WX8944,WX8943,WX8945,WX8949,WX8951,WX8950,WX8952,
    WX8956,WX8958,WX8957,WX8959,WX8963,WX8965,WX8964,WX8966,WX8970,WX8972,
    WX8971,WX8973,WX8977,WX8979,WX8978,WX8980,WX8984,WX8986,WX8985,WX8987,
    WX8988,WX9021,WX9088,WX10054,WX9092,WX10055,WX9096,WX9098,WX9089,WX9099,
    WX9102,WX9106,WX9110,WX9112,WX9103,WX9113,WX9116,WX9120,WX9124,WX9126,
    WX9117,WX9127,WX9130,WX9134,WX9138,WX9140,WX9131,WX9141,WX9144,WX9148,
    WX9152,WX9154,WX9145,WX9155,WX9158,WX9162,WX9166,WX9168,WX9159,WX9169,
    WX9172,WX9176,WX9180,WX9182,WX9173,WX9183,WX9186,WX9190,WX9194,WX9196,
    WX9187,WX9197,WX9200,WX9204,WX9208,WX9210,WX9201,WX9211,WX9214,WX9218,
    WX9222,WX9224,WX9215,WX9225,WX9228,WX9232,WX9236,WX9238,WX9229,WX9239,
    WX9242,WX9246,WX9250,WX9252,WX9243,WX9253,WX9256,WX9260,WX9264,WX9266,
    WX9257,WX9267,WX9270,WX9274,WX9278,WX9280,WX9271,WX9281,WX9284,WX9288,
    WX9292,WX9294,WX9285,WX9295,WX9298,WX9302,WX9306,WX9308,WX9299,WX9309,
    WX9312,WX9316,WX9320,WX9322,WX9313,WX9323,WX9326,WX9330,WX9334,WX9336,
    WX9327,WX9337,WX9340,WX9344,WX9348,WX9350,WX9341,WX9351,WX9354,WX9358,
    WX9362,WX9364,WX9355,WX9365,WX9368,WX9372,WX9376,WX9378,WX9369,WX9379,
    WX9382,WX9386,WX9390,WX9392,WX9383,WX9393,WX9396,WX9400,WX9404,WX9406,
    WX9397,WX9407,WX9410,WX9414,WX9418,WX9420,WX9411,WX9421,WX9424,WX9428,
    WX9432,WX9434,WX9425,WX9435,WX9438,WX9442,WX9446,WX9448,WX9439,WX9449,
    WX9452,WX9456,WX9460,WX9462,WX9453,WX9463,WX9466,WX9470,WX9474,WX9476,
    WX9467,WX9477,WX9480,WX9484,WX9488,WX9490,WX9481,WX9491,WX9494,WX9498,
    WX9502,WX9504,WX9495,WX9505,WX9508,WX9512,WX9516,WX9518,WX9509,WX9519,
    WX9522,WX9526,WX9530,WX9532,WX9523,WX9533,WX9534,WX9599,WX10016,WX9600,
    WX10018,WX9601,WX10020,WX9602,WX10022,WX9603,WX10024,WX9604,WX10026,WX9605,
    WX10028,WX9606,WX10030,WX9607,WX10032,WX9608,WX10034,WX9609,WX10036,WX9610,
    WX10038,WX9611,WX10040,WX9612,WX10042,WX9613,WX10044,WX9614,WX10046,WX9615,
    WX9984,WX9616,WX9986,WX9617,WX9988,WX9618,WX9990,WX9619,WX9992,WX9620,
    WX9994,WX9621,WX9996,WX9622,WX9998,WX9623,WX10000,WX9624,WX10002,WX9625,
    WX10004,WX9626,WX10006,WX9627,WX10008,WX9628,WX10010,WX9629,WX10012,WX9630,
    WX10014,WX9631,WX9632,WX9633,WX9634,WX9635,WX9636,WX9637,WX9638,WX9639,
    WX9640,WX9641,WX9642,WX9643,WX9644,WX9645,WX9646,WX9647,WX9648,WX9649,
    WX9650,WX9651,WX9652,WX9653,WX9654,WX9655,WX9656,WX9657,WX9658,WX9659,
    WX9660,WX9661,WX9662,WX9663,WX9664,WX9665,WX9666,WX9667,WX9668,WX9669,
    WX9670,WX9671,WX9672,WX9673,WX9674,WX9675,WX9676,WX9677,WX9678,WX9679,
    WX9680,WX9681,WX9682,WX9683,WX9684,WX9685,WX9686,WX9687,WX9688,WX9689,
    WX9690,WX9691,WX9692,WX9693,WX9694,WX9983,WX9967,WX9985,WX9968,WX9987,
    WX9969,WX9989,WX9970,WX9991,WX9971,WX9993,WX9972,WX9995,WX9973,WX9997,
    WX9974,WX9999,WX9975,WX10001,WX9976,WX10003,WX9977,WX10005,WX9978,WX10007,
    WX9979,WX10009,WX9980,WX10011,WX9981,WX10013,WX9982,WX10015,WX9951,WX10017,
    WX9952,WX10019,WX9953,WX10021,WX9954,WX10023,WX9955,WX10025,WX9956,WX10027,
    WX9957,WX10029,WX9958,WX10031,WX9959,WX10033,WX9960,WX10035,WX9961,WX10037,
    WX9962,WX10039,WX9963,WX10041,WX9964,WX10043,WX9965,WX10045,WX9966,WX10047,
    WX10048,WX10049,WX10050,WX10051,WX10052,WX10053,WX10056,WX10060,WX10062,
    WX10061,WX10063,WX10067,WX10069,WX10068,WX10070,WX10074,WX10076,WX10075,
    WX10077,WX10081,WX10083,WX10082,WX10084,WX10088,WX10090,WX10089,WX10091,
    WX10095,WX10097,WX10096,WX10098,WX10102,WX10104,WX10103,WX10105,WX10109,
    WX10111,WX10110,WX10112,WX10116,WX10118,WX10117,WX10119,WX10123,WX10125,
    WX10124,WX10126,WX10130,WX10132,WX10131,WX10133,WX10137,WX10139,WX10138,
    WX10140,WX10144,WX10146,WX10145,WX10147,WX10151,WX10153,WX10152,WX10154,
    WX10158,WX10160,WX10159,WX10161,WX10165,WX10167,WX10166,WX10168,WX10172,
    WX10174,WX10173,WX10175,WX10179,WX10181,WX10180,WX10182,WX10186,WX10188,
    WX10187,WX10189,WX10193,WX10195,WX10194,WX10196,WX10200,WX10202,WX10201,
    WX10203,WX10207,WX10209,WX10208,WX10210,WX10214,WX10216,WX10215,WX10217,
    WX10221,WX10223,WX10222,WX10224,WX10228,WX10230,WX10229,WX10231,WX10235,
    WX10237,WX10236,WX10238,WX10242,WX10244,WX10243,WX10245,WX10249,WX10251,
    WX10250,WX10252,WX10256,WX10258,WX10257,WX10259,WX10263,WX10265,WX10264,
    WX10266,WX10270,WX10272,WX10271,WX10273,WX10277,WX10279,WX10278,WX10280,
    WX10281,WX10314,WX10381,WX11347,WX10385,WX11348,WX10389,WX10391,WX10382,
    WX10392,WX10395,WX10399,WX10403,WX10405,WX10396,WX10406,WX10409,WX10413,
    WX10417,WX10419,WX10410,WX10420,WX10423,WX10427,WX10431,WX10433,WX10424,
    WX10434,WX10437,WX10441,WX10445,WX10447,WX10438,WX10448,WX10451,WX10455,
    WX10459,WX10461,WX10452,WX10462,WX10465,WX10469,WX10473,WX10475,WX10466,
    WX10476,WX10479,WX10483,WX10487,WX10489,WX10480,WX10490,WX10493,WX10497,
    WX10501,WX10503,WX10494,WX10504,WX10507,WX10511,WX10515,WX10517,WX10508,
    WX10518,WX10521,WX10525,WX10529,WX10531,WX10522,WX10532,WX10535,WX10539,
    WX10543,WX10545,WX10536,WX10546,WX10549,WX10553,WX10557,WX10559,WX10550,
    WX10560,WX10563,WX10567,WX10571,WX10573,WX10564,WX10574,WX10577,WX10581,
    WX10585,WX10587,WX10578,WX10588,WX10591,WX10595,WX10599,WX10601,WX10592,
    WX10602,WX10605,WX10609,WX10613,WX10615,WX10606,WX10616,WX10619,WX10623,
    WX10627,WX10629,WX10620,WX10630,WX10633,WX10637,WX10641,WX10643,WX10634,
    WX10644,WX10647,WX10651,WX10655,WX10657,WX10648,WX10658,WX10661,WX10665,
    WX10669,WX10671,WX10662,WX10672,WX10675,WX10679,WX10683,WX10685,WX10676,
    WX10686,WX10689,WX10693,WX10697,WX10699,WX10690,WX10700,WX10703,WX10707,
    WX10711,WX10713,WX10704,WX10714,WX10717,WX10721,WX10725,WX10727,WX10718,
    WX10728,WX10731,WX10735,WX10739,WX10741,WX10732,WX10742,WX10745,WX10749,
    WX10753,WX10755,WX10746,WX10756,WX10759,WX10763,WX10767,WX10769,WX10760,
    WX10770,WX10773,WX10777,WX10781,WX10783,WX10774,WX10784,WX10787,WX10791,
    WX10795,WX10797,WX10788,WX10798,WX10801,WX10805,WX10809,WX10811,WX10802,
    WX10812,WX10815,WX10819,WX10823,WX10825,WX10816,WX10826,WX10827,WX10892,
    WX11309,WX10893,WX11311,WX10894,WX11313,WX10895,WX11315,WX10896,WX11317,
    WX10897,WX11319,WX10898,WX11321,WX10899,WX11323,WX10900,WX11325,WX10901,
    WX11327,WX10902,WX11329,WX10903,WX11331,WX10904,WX11333,WX10905,WX11335,
    WX10906,WX11337,WX10907,WX11339,WX10908,WX11277,WX10909,WX11279,WX10910,
    WX11281,WX10911,WX11283,WX10912,WX11285,WX10913,WX11287,WX10914,WX11289,
    WX10915,WX11291,WX10916,WX11293,WX10917,WX11295,WX10918,WX11297,WX10919,
    WX11299,WX10920,WX11301,WX10921,WX11303,WX10922,WX11305,WX10923,WX11307,
    WX10924,WX10925,WX10926,WX10927,WX10928,WX10929,WX10930,WX10931,WX10932,
    WX10933,WX10934,WX10935,WX10936,WX10937,WX10938,WX10939,WX10940,WX10941,
    WX10942,WX10943,WX10944,WX10945,WX10946,WX10947,WX10948,WX10949,WX10950,
    WX10951,WX10952,WX10953,WX10954,WX10955,WX10956,WX10957,WX10958,WX10959,
    WX10960,WX10961,WX10962,WX10963,WX10964,WX10965,WX10966,WX10967,WX10968,
    WX10969,WX10970,WX10971,WX10972,WX10973,WX10974,WX10975,WX10976,WX10977,
    WX10978,WX10979,WX10980,WX10981,WX10982,WX10983,WX10984,WX10985,WX10986,
    WX10987,WX11276,WX11260,WX11278,WX11261,WX11280,WX11262,WX11282,WX11263,
    WX11284,WX11264,WX11286,WX11265,WX11288,WX11266,WX11290,WX11267,WX11292,
    WX11268,WX11294,WX11269,WX11296,WX11270,WX11298,WX11271,WX11300,WX11272,
    WX11302,WX11273,WX11304,WX11274,WX11306,WX11275,WX11308,WX11244,WX11310,
    WX11245,WX11312,WX11246,WX11314,WX11247,WX11316,WX11248,WX11318,WX11249,
    WX11320,WX11250,WX11322,WX11251,WX11324,WX11252,WX11326,WX11253,WX11328,
    WX11254,WX11330,WX11255,WX11332,WX11256,WX11334,WX11257,WX11336,WX11258,
    WX11338,WX11259,WX11340,WX11341,WX11342,WX11343,WX11344,WX11345,WX11346,
    WX11349,WX11353,WX11355,WX11354,WX11356,WX11360,WX11362,WX11361,WX11363,
    WX11367,WX11369,WX11368,WX11370,WX11374,WX11376,WX11375,WX11377,WX11381,
    WX11383,WX11382,WX11384,WX11388,WX11390,WX11389,WX11391,WX11395,WX11397,
    WX11396,WX11398,WX11402,WX11404,WX11403,WX11405,WX11409,WX11411,WX11410,
    WX11412,WX11416,WX11418,WX11417,WX11419,WX11423,WX11425,WX11424,WX11426,
    WX11430,WX11432,WX11431,WX11433,WX11437,WX11439,WX11438,WX11440,WX11444,
    WX11446,WX11445,WX11447,WX11451,WX11453,WX11452,WX11454,WX11458,WX11460,
    WX11459,WX11461,WX11465,WX11467,WX11466,WX11468,WX11472,WX11474,WX11473,
    WX11475,WX11479,WX11481,WX11480,WX11482,WX11486,WX11488,WX11487,WX11489,
    WX11493,WX11495,WX11494,WX11496,WX11500,WX11502,WX11501,WX11503,WX11507,
    WX11509,WX11508,WX11510,WX11514,WX11516,WX11515,WX11517,WX11521,WX11523,
    WX11522,WX11524,WX11528,WX11530,WX11529,WX11531,WX11535,WX11537,WX11536,
    WX11538,WX11542,WX11544,WX11543,WX11545,WX11549,WX11551,WX11550,WX11552,
    WX11556,WX11558,WX11557,WX11559,WX11563,WX11565,WX11564,WX11566,WX11570,
    WX11572,WX11571,WX11573,WX11574,WX11607,WX35,WX46,WX36,WX42,WX39,WX40,WX43,
    WX44,WX49,WX60,WX50,WX56,WX53,WX54,WX57,WX58,WX63,WX74,WX64,WX70,WX67,WX68,
    WX71,WX72,WX77,WX88,WX78,WX84,WX81,WX82,WX85,WX86,WX91,WX102,WX92,WX98,
    WX95,WX96,WX99,WX100,WX105,WX116,WX106,WX112,WX109,WX110,WX113,WX114,WX119,
    WX130,WX120,WX126,WX123,WX124,WX127,WX128,WX133,WX144,WX134,WX140,WX137,
    WX138,WX141,WX142,WX147,WX158,WX148,WX154,WX151,WX152,WX155,WX156,WX161,
    WX172,WX162,WX168,WX165,WX166,WX169,WX170,WX175,WX186,WX176,WX182,WX179,
    WX180,WX183,WX184,WX189,WX200,WX190,WX196,WX193,WX194,WX197,WX198,WX203,
    WX214,WX204,WX210,WX207,WX208,WX211,WX212,WX217,WX228,WX218,WX224,WX221,
    WX222,WX225,WX226,WX231,WX242,WX232,WX238,WX235,WX236,WX239,WX240,WX245,
    WX256,WX246,WX252,WX249,WX250,WX253,WX254,WX259,WX270,WX260,WX266,WX263,
    WX264,WX267,WX268,WX273,WX284,WX274,WX280,WX277,WX278,WX281,WX282,WX287,
    WX298,WX288,WX294,WX291,WX292,WX295,WX296,WX301,WX312,WX302,WX308,WX305,
    WX306,WX309,WX310,WX315,WX326,WX316,WX322,WX319,WX320,WX323,WX324,WX329,
    WX340,WX330,WX336,WX333,WX334,WX337,WX338,WX343,WX354,WX344,WX350,WX347,
    WX348,WX351,WX352,WX357,WX368,WX358,WX364,WX361,WX362,WX365,WX366,WX371,
    WX382,WX372,WX378,WX375,WX376,WX379,WX380,WX385,WX396,WX386,WX392,WX389,
    WX390,WX393,WX394,WX399,WX410,WX400,WX406,WX403,WX404,WX407,WX408,WX413,
    WX424,WX414,WX420,WX417,WX418,WX421,WX422,WX427,WX438,WX428,WX434,WX431,
    WX432,WX435,WX436,WX441,WX452,WX442,WX448,WX445,WX446,WX449,WX450,WX455,
    WX466,WX456,WX462,WX459,WX460,WX463,WX464,WX469,WX480,WX470,WX476,WX473,
    WX474,WX477,WX478,WX1007,WX1006,WX1008,WX1014,WX1013,WX1015,WX1021,WX1020,
    WX1022,WX1028,WX1027,WX1029,WX1035,WX1034,WX1036,WX1042,WX1041,WX1043,
    WX1049,WX1048,WX1050,WX1056,WX1055,WX1057,WX1063,WX1062,WX1064,WX1070,
    WX1069,WX1071,WX1077,WX1076,WX1078,WX1084,WX1083,WX1085,WX1091,WX1090,
    WX1092,WX1098,WX1097,WX1099,WX1105,WX1104,WX1106,WX1112,WX1111,WX1113,
    WX1119,WX1118,WX1120,WX1126,WX1125,WX1127,WX1133,WX1132,WX1134,WX1140,
    WX1139,WX1141,WX1147,WX1146,WX1148,WX1154,WX1153,WX1155,WX1161,WX1160,
    WX1162,WX1168,WX1167,WX1169,WX1175,WX1174,WX1176,WX1182,WX1181,WX1183,
    WX1189,WX1188,WX1190,WX1196,WX1195,WX1197,WX1203,WX1202,WX1204,WX1210,
    WX1209,WX1211,WX1217,WX1216,WX1218,WX1224,WX1223,WX1225,WX1234,WX1262,
    WX1261,WX1260,WX1233,WX1259,WX1258,WX1257,WX1256,WX1255,WX1254,WX1232,
    WX1253,WX1252,WX1251,WX1250,WX1231,WX1249,WX1248,WX1247,WX1246,WX1245,
    WX1244,WX1243,WX1242,WX1241,WX1240,WX1239,WX1238,WX1237,WX1236,WX1235,
    WX1328,WX1339,WX1329,WX1335,WX1332,WX1333,WX1336,WX1337,WX1342,WX1353,
    WX1343,WX1349,WX1346,WX1347,WX1350,WX1351,WX1356,WX1367,WX1357,WX1363,
    WX1360,WX1361,WX1364,WX1365,WX1370,WX1381,WX1371,WX1377,WX1374,WX1375,
    WX1378,WX1379,WX1384,WX1395,WX1385,WX1391,WX1388,WX1389,WX1392,WX1393,
    WX1398,WX1409,WX1399,WX1405,WX1402,WX1403,WX1406,WX1407,WX1412,WX1423,
    WX1413,WX1419,WX1416,WX1417,WX1420,WX1421,WX1426,WX1437,WX1427,WX1433,
    WX1430,WX1431,WX1434,WX1435,WX1440,WX1451,WX1441,WX1447,WX1444,WX1445,
    WX1448,WX1449,WX1454,WX1465,WX1455,WX1461,WX1458,WX1459,WX1462,WX1463,
    WX1468,WX1479,WX1469,WX1475,WX1472,WX1473,WX1476,WX1477,WX1482,WX1493,
    WX1483,WX1489,WX1486,WX1487,WX1490,WX1491,WX1496,WX1507,WX1497,WX1503,
    WX1500,WX1501,WX1504,WX1505,WX1510,WX1521,WX1511,WX1517,WX1514,WX1515,
    WX1518,WX1519,WX1524,WX1535,WX1525,WX1531,WX1528,WX1529,WX1532,WX1533,
    WX1538,WX1549,WX1539,WX1545,WX1542,WX1543,WX1546,WX1547,WX1552,WX1563,
    WX1553,WX1559,WX1556,WX1557,WX1560,WX1561,WX1566,WX1577,WX1567,WX1573,
    WX1570,WX1571,WX1574,WX1575,WX1580,WX1591,WX1581,WX1587,WX1584,WX1585,
    WX1588,WX1589,WX1594,WX1605,WX1595,WX1601,WX1598,WX1599,WX1602,WX1603,
    WX1608,WX1619,WX1609,WX1615,WX1612,WX1613,WX1616,WX1617,WX1622,WX1633,
    WX1623,WX1629,WX1626,WX1627,WX1630,WX1631,WX1636,WX1647,WX1637,WX1643,
    WX1640,WX1641,WX1644,WX1645,WX1650,WX1661,WX1651,WX1657,WX1654,WX1655,
    WX1658,WX1659,WX1664,WX1675,WX1665,WX1671,WX1668,WX1669,WX1672,WX1673,
    WX1678,WX1689,WX1679,WX1685,WX1682,WX1683,WX1686,WX1687,WX1692,WX1703,
    WX1693,WX1699,WX1696,WX1697,WX1700,WX1701,WX1706,WX1717,WX1707,WX1713,
    WX1710,WX1711,WX1714,WX1715,WX1720,WX1731,WX1721,WX1727,WX1724,WX1725,
    WX1728,WX1729,WX1734,WX1745,WX1735,WX1741,WX1738,WX1739,WX1742,WX1743,
    WX1748,WX1759,WX1749,WX1755,WX1752,WX1753,WX1756,WX1757,WX1762,WX1773,
    WX1763,WX1769,WX1766,WX1767,WX1770,WX1771,WX2300,WX2299,WX2301,WX2307,
    WX2306,WX2308,WX2314,WX2313,WX2315,WX2321,WX2320,WX2322,WX2328,WX2327,
    WX2329,WX2335,WX2334,WX2336,WX2342,WX2341,WX2343,WX2349,WX2348,WX2350,
    WX2356,WX2355,WX2357,WX2363,WX2362,WX2364,WX2370,WX2369,WX2371,WX2377,
    WX2376,WX2378,WX2384,WX2383,WX2385,WX2391,WX2390,WX2392,WX2398,WX2397,
    WX2399,WX2405,WX2404,WX2406,WX2412,WX2411,WX2413,WX2419,WX2418,WX2420,
    WX2426,WX2425,WX2427,WX2433,WX2432,WX2434,WX2440,WX2439,WX2441,WX2447,
    WX2446,WX2448,WX2454,WX2453,WX2455,WX2461,WX2460,WX2462,WX2468,WX2467,
    WX2469,WX2475,WX2474,WX2476,WX2482,WX2481,WX2483,WX2489,WX2488,WX2490,
    WX2496,WX2495,WX2497,WX2503,WX2502,WX2504,WX2510,WX2509,WX2511,WX2517,
    WX2516,WX2518,WX2527,WX2555,WX2554,WX2553,WX2526,WX2552,WX2551,WX2550,
    WX2549,WX2548,WX2547,WX2525,WX2546,WX2545,WX2544,WX2543,WX2524,WX2542,
    WX2541,WX2540,WX2539,WX2538,WX2537,WX2536,WX2535,WX2534,WX2533,WX2532,
    WX2531,WX2530,WX2529,WX2528,WX2621,WX2632,WX2622,WX2628,WX2625,WX2626,
    WX2629,WX2630,WX2635,WX2646,WX2636,WX2642,WX2639,WX2640,WX2643,WX2644,
    WX2649,WX2660,WX2650,WX2656,WX2653,WX2654,WX2657,WX2658,WX2663,WX2674,
    WX2664,WX2670,WX2667,WX2668,WX2671,WX2672,WX2677,WX2688,WX2678,WX2684,
    WX2681,WX2682,WX2685,WX2686,WX2691,WX2702,WX2692,WX2698,WX2695,WX2696,
    WX2699,WX2700,WX2705,WX2716,WX2706,WX2712,WX2709,WX2710,WX2713,WX2714,
    WX2719,WX2730,WX2720,WX2726,WX2723,WX2724,WX2727,WX2728,WX2733,WX2744,
    WX2734,WX2740,WX2737,WX2738,WX2741,WX2742,WX2747,WX2758,WX2748,WX2754,
    WX2751,WX2752,WX2755,WX2756,WX2761,WX2772,WX2762,WX2768,WX2765,WX2766,
    WX2769,WX2770,WX2775,WX2786,WX2776,WX2782,WX2779,WX2780,WX2783,WX2784,
    WX2789,WX2800,WX2790,WX2796,WX2793,WX2794,WX2797,WX2798,WX2803,WX2814,
    WX2804,WX2810,WX2807,WX2808,WX2811,WX2812,WX2817,WX2828,WX2818,WX2824,
    WX2821,WX2822,WX2825,WX2826,WX2831,WX2842,WX2832,WX2838,WX2835,WX2836,
    WX2839,WX2840,WX2845,WX2856,WX2846,WX2852,WX2849,WX2850,WX2853,WX2854,
    WX2859,WX2870,WX2860,WX2866,WX2863,WX2864,WX2867,WX2868,WX2873,WX2884,
    WX2874,WX2880,WX2877,WX2878,WX2881,WX2882,WX2887,WX2898,WX2888,WX2894,
    WX2891,WX2892,WX2895,WX2896,WX2901,WX2912,WX2902,WX2908,WX2905,WX2906,
    WX2909,WX2910,WX2915,WX2926,WX2916,WX2922,WX2919,WX2920,WX2923,WX2924,
    WX2929,WX2940,WX2930,WX2936,WX2933,WX2934,WX2937,WX2938,WX2943,WX2954,
    WX2944,WX2950,WX2947,WX2948,WX2951,WX2952,WX2957,WX2968,WX2958,WX2964,
    WX2961,WX2962,WX2965,WX2966,WX2971,WX2982,WX2972,WX2978,WX2975,WX2976,
    WX2979,WX2980,WX2985,WX2996,WX2986,WX2992,WX2989,WX2990,WX2993,WX2994,
    WX2999,WX3010,WX3000,WX3006,WX3003,WX3004,WX3007,WX3008,WX3013,WX3024,
    WX3014,WX3020,WX3017,WX3018,WX3021,WX3022,WX3027,WX3038,WX3028,WX3034,
    WX3031,WX3032,WX3035,WX3036,WX3041,WX3052,WX3042,WX3048,WX3045,WX3046,
    WX3049,WX3050,WX3055,WX3066,WX3056,WX3062,WX3059,WX3060,WX3063,WX3064,
    WX3593,WX3592,WX3594,WX3600,WX3599,WX3601,WX3607,WX3606,WX3608,WX3614,
    WX3613,WX3615,WX3621,WX3620,WX3622,WX3628,WX3627,WX3629,WX3635,WX3634,
    WX3636,WX3642,WX3641,WX3643,WX3649,WX3648,WX3650,WX3656,WX3655,WX3657,
    WX3663,WX3662,WX3664,WX3670,WX3669,WX3671,WX3677,WX3676,WX3678,WX3684,
    WX3683,WX3685,WX3691,WX3690,WX3692,WX3698,WX3697,WX3699,WX3705,WX3704,
    WX3706,WX3712,WX3711,WX3713,WX3719,WX3718,WX3720,WX3726,WX3725,WX3727,
    WX3733,WX3732,WX3734,WX3740,WX3739,WX3741,WX3747,WX3746,WX3748,WX3754,
    WX3753,WX3755,WX3761,WX3760,WX3762,WX3768,WX3767,WX3769,WX3775,WX3774,
    WX3776,WX3782,WX3781,WX3783,WX3789,WX3788,WX3790,WX3796,WX3795,WX3797,
    WX3803,WX3802,WX3804,WX3810,WX3809,WX3811,WX3820,WX3848,WX3847,WX3846,
    WX3819,WX3845,WX3844,WX3843,WX3842,WX3841,WX3840,WX3818,WX3839,WX3838,
    WX3837,WX3836,WX3817,WX3835,WX3834,WX3833,WX3832,WX3831,WX3830,WX3829,
    WX3828,WX3827,WX3826,WX3825,WX3824,WX3823,WX3822,WX3821,WX3914,WX3925,
    WX3915,WX3921,WX3918,WX3919,WX3922,WX3923,WX3928,WX3939,WX3929,WX3935,
    WX3932,WX3933,WX3936,WX3937,WX3942,WX3953,WX3943,WX3949,WX3946,WX3947,
    WX3950,WX3951,WX3956,WX3967,WX3957,WX3963,WX3960,WX3961,WX3964,WX3965,
    WX3970,WX3981,WX3971,WX3977,WX3974,WX3975,WX3978,WX3979,WX3984,WX3995,
    WX3985,WX3991,WX3988,WX3989,WX3992,WX3993,WX3998,WX4009,WX3999,WX4005,
    WX4002,WX4003,WX4006,WX4007,WX4012,WX4023,WX4013,WX4019,WX4016,WX4017,
    WX4020,WX4021,WX4026,WX4037,WX4027,WX4033,WX4030,WX4031,WX4034,WX4035,
    WX4040,WX4051,WX4041,WX4047,WX4044,WX4045,WX4048,WX4049,WX4054,WX4065,
    WX4055,WX4061,WX4058,WX4059,WX4062,WX4063,WX4068,WX4079,WX4069,WX4075,
    WX4072,WX4073,WX4076,WX4077,WX4082,WX4093,WX4083,WX4089,WX4086,WX4087,
    WX4090,WX4091,WX4096,WX4107,WX4097,WX4103,WX4100,WX4101,WX4104,WX4105,
    WX4110,WX4121,WX4111,WX4117,WX4114,WX4115,WX4118,WX4119,WX4124,WX4135,
    WX4125,WX4131,WX4128,WX4129,WX4132,WX4133,WX4138,WX4149,WX4139,WX4145,
    WX4142,WX4143,WX4146,WX4147,WX4152,WX4163,WX4153,WX4159,WX4156,WX4157,
    WX4160,WX4161,WX4166,WX4177,WX4167,WX4173,WX4170,WX4171,WX4174,WX4175,
    WX4180,WX4191,WX4181,WX4187,WX4184,WX4185,WX4188,WX4189,WX4194,WX4205,
    WX4195,WX4201,WX4198,WX4199,WX4202,WX4203,WX4208,WX4219,WX4209,WX4215,
    WX4212,WX4213,WX4216,WX4217,WX4222,WX4233,WX4223,WX4229,WX4226,WX4227,
    WX4230,WX4231,WX4236,WX4247,WX4237,WX4243,WX4240,WX4241,WX4244,WX4245,
    WX4250,WX4261,WX4251,WX4257,WX4254,WX4255,WX4258,WX4259,WX4264,WX4275,
    WX4265,WX4271,WX4268,WX4269,WX4272,WX4273,WX4278,WX4289,WX4279,WX4285,
    WX4282,WX4283,WX4286,WX4287,WX4292,WX4303,WX4293,WX4299,WX4296,WX4297,
    WX4300,WX4301,WX4306,WX4317,WX4307,WX4313,WX4310,WX4311,WX4314,WX4315,
    WX4320,WX4331,WX4321,WX4327,WX4324,WX4325,WX4328,WX4329,WX4334,WX4345,
    WX4335,WX4341,WX4338,WX4339,WX4342,WX4343,WX4348,WX4359,WX4349,WX4355,
    WX4352,WX4353,WX4356,WX4357,WX4886,WX4885,WX4887,WX4893,WX4892,WX4894,
    WX4900,WX4899,WX4901,WX4907,WX4906,WX4908,WX4914,WX4913,WX4915,WX4921,
    WX4920,WX4922,WX4928,WX4927,WX4929,WX4935,WX4934,WX4936,WX4942,WX4941,
    WX4943,WX4949,WX4948,WX4950,WX4956,WX4955,WX4957,WX4963,WX4962,WX4964,
    WX4970,WX4969,WX4971,WX4977,WX4976,WX4978,WX4984,WX4983,WX4985,WX4991,
    WX4990,WX4992,WX4998,WX4997,WX4999,WX5005,WX5004,WX5006,WX5012,WX5011,
    WX5013,WX5019,WX5018,WX5020,WX5026,WX5025,WX5027,WX5033,WX5032,WX5034,
    WX5040,WX5039,WX5041,WX5047,WX5046,WX5048,WX5054,WX5053,WX5055,WX5061,
    WX5060,WX5062,WX5068,WX5067,WX5069,WX5075,WX5074,WX5076,WX5082,WX5081,
    WX5083,WX5089,WX5088,WX5090,WX5096,WX5095,WX5097,WX5103,WX5102,WX5104,
    WX5113,WX5141,WX5140,WX5139,WX5112,WX5138,WX5137,WX5136,WX5135,WX5134,
    WX5133,WX5111,WX5132,WX5131,WX5130,WX5129,WX5110,WX5128,WX5127,WX5126,
    WX5125,WX5124,WX5123,WX5122,WX5121,WX5120,WX5119,WX5118,WX5117,WX5116,
    WX5115,WX5114,WX5207,WX5218,WX5208,WX5214,WX5211,WX5212,WX5215,WX5216,
    WX5221,WX5232,WX5222,WX5228,WX5225,WX5226,WX5229,WX5230,WX5235,WX5246,
    WX5236,WX5242,WX5239,WX5240,WX5243,WX5244,WX5249,WX5260,WX5250,WX5256,
    WX5253,WX5254,WX5257,WX5258,WX5263,WX5274,WX5264,WX5270,WX5267,WX5268,
    WX5271,WX5272,WX5277,WX5288,WX5278,WX5284,WX5281,WX5282,WX5285,WX5286,
    WX5291,WX5302,WX5292,WX5298,WX5295,WX5296,WX5299,WX5300,WX5305,WX5316,
    WX5306,WX5312,WX5309,WX5310,WX5313,WX5314,WX5319,WX5330,WX5320,WX5326,
    WX5323,WX5324,WX5327,WX5328,WX5333,WX5344,WX5334,WX5340,WX5337,WX5338,
    WX5341,WX5342,WX5347,WX5358,WX5348,WX5354,WX5351,WX5352,WX5355,WX5356,
    WX5361,WX5372,WX5362,WX5368,WX5365,WX5366,WX5369,WX5370,WX5375,WX5386,
    WX5376,WX5382,WX5379,WX5380,WX5383,WX5384,WX5389,WX5400,WX5390,WX5396,
    WX5393,WX5394,WX5397,WX5398,WX5403,WX5414,WX5404,WX5410,WX5407,WX5408,
    WX5411,WX5412,WX5417,WX5428,WX5418,WX5424,WX5421,WX5422,WX5425,WX5426,
    WX5431,WX5442,WX5432,WX5438,WX5435,WX5436,WX5439,WX5440,WX5445,WX5456,
    WX5446,WX5452,WX5449,WX5450,WX5453,WX5454,WX5459,WX5470,WX5460,WX5466,
    WX5463,WX5464,WX5467,WX5468,WX5473,WX5484,WX5474,WX5480,WX5477,WX5478,
    WX5481,WX5482,WX5487,WX5498,WX5488,WX5494,WX5491,WX5492,WX5495,WX5496,
    WX5501,WX5512,WX5502,WX5508,WX5505,WX5506,WX5509,WX5510,WX5515,WX5526,
    WX5516,WX5522,WX5519,WX5520,WX5523,WX5524,WX5529,WX5540,WX5530,WX5536,
    WX5533,WX5534,WX5537,WX5538,WX5543,WX5554,WX5544,WX5550,WX5547,WX5548,
    WX5551,WX5552,WX5557,WX5568,WX5558,WX5564,WX5561,WX5562,WX5565,WX5566,
    WX5571,WX5582,WX5572,WX5578,WX5575,WX5576,WX5579,WX5580,WX5585,WX5596,
    WX5586,WX5592,WX5589,WX5590,WX5593,WX5594,WX5599,WX5610,WX5600,WX5606,
    WX5603,WX5604,WX5607,WX5608,WX5613,WX5624,WX5614,WX5620,WX5617,WX5618,
    WX5621,WX5622,WX5627,WX5638,WX5628,WX5634,WX5631,WX5632,WX5635,WX5636,
    WX5641,WX5652,WX5642,WX5648,WX5645,WX5646,WX5649,WX5650,WX6179,WX6178,
    WX6180,WX6186,WX6185,WX6187,WX6193,WX6192,WX6194,WX6200,WX6199,WX6201,
    WX6207,WX6206,WX6208,WX6214,WX6213,WX6215,WX6221,WX6220,WX6222,WX6228,
    WX6227,WX6229,WX6235,WX6234,WX6236,WX6242,WX6241,WX6243,WX6249,WX6248,
    WX6250,WX6256,WX6255,WX6257,WX6263,WX6262,WX6264,WX6270,WX6269,WX6271,
    WX6277,WX6276,WX6278,WX6284,WX6283,WX6285,WX6291,WX6290,WX6292,WX6298,
    WX6297,WX6299,WX6305,WX6304,WX6306,WX6312,WX6311,WX6313,WX6319,WX6318,
    WX6320,WX6326,WX6325,WX6327,WX6333,WX6332,WX6334,WX6340,WX6339,WX6341,
    WX6347,WX6346,WX6348,WX6354,WX6353,WX6355,WX6361,WX6360,WX6362,WX6368,
    WX6367,WX6369,WX6375,WX6374,WX6376,WX6382,WX6381,WX6383,WX6389,WX6388,
    WX6390,WX6396,WX6395,WX6397,WX6406,WX6434,WX6433,WX6432,WX6405,WX6431,
    WX6430,WX6429,WX6428,WX6427,WX6426,WX6404,WX6425,WX6424,WX6423,WX6422,
    WX6403,WX6421,WX6420,WX6419,WX6418,WX6417,WX6416,WX6415,WX6414,WX6413,
    WX6412,WX6411,WX6410,WX6409,WX6408,WX6407,WX6500,WX6511,WX6501,WX6507,
    WX6504,WX6505,WX6508,WX6509,WX6514,WX6525,WX6515,WX6521,WX6518,WX6519,
    WX6522,WX6523,WX6528,WX6539,WX6529,WX6535,WX6532,WX6533,WX6536,WX6537,
    WX6542,WX6553,WX6543,WX6549,WX6546,WX6547,WX6550,WX6551,WX6556,WX6567,
    WX6557,WX6563,WX6560,WX6561,WX6564,WX6565,WX6570,WX6581,WX6571,WX6577,
    WX6574,WX6575,WX6578,WX6579,WX6584,WX6595,WX6585,WX6591,WX6588,WX6589,
    WX6592,WX6593,WX6598,WX6609,WX6599,WX6605,WX6602,WX6603,WX6606,WX6607,
    WX6612,WX6623,WX6613,WX6619,WX6616,WX6617,WX6620,WX6621,WX6626,WX6637,
    WX6627,WX6633,WX6630,WX6631,WX6634,WX6635,WX6640,WX6651,WX6641,WX6647,
    WX6644,WX6645,WX6648,WX6649,WX6654,WX6665,WX6655,WX6661,WX6658,WX6659,
    WX6662,WX6663,WX6668,WX6679,WX6669,WX6675,WX6672,WX6673,WX6676,WX6677,
    WX6682,WX6693,WX6683,WX6689,WX6686,WX6687,WX6690,WX6691,WX6696,WX6707,
    WX6697,WX6703,WX6700,WX6701,WX6704,WX6705,WX6710,WX6721,WX6711,WX6717,
    WX6714,WX6715,WX6718,WX6719,WX6724,WX6735,WX6725,WX6731,WX6728,WX6729,
    WX6732,WX6733,WX6738,WX6749,WX6739,WX6745,WX6742,WX6743,WX6746,WX6747,
    WX6752,WX6763,WX6753,WX6759,WX6756,WX6757,WX6760,WX6761,WX6766,WX6777,
    WX6767,WX6773,WX6770,WX6771,WX6774,WX6775,WX6780,WX6791,WX6781,WX6787,
    WX6784,WX6785,WX6788,WX6789,WX6794,WX6805,WX6795,WX6801,WX6798,WX6799,
    WX6802,WX6803,WX6808,WX6819,WX6809,WX6815,WX6812,WX6813,WX6816,WX6817,
    WX6822,WX6833,WX6823,WX6829,WX6826,WX6827,WX6830,WX6831,WX6836,WX6847,
    WX6837,WX6843,WX6840,WX6841,WX6844,WX6845,WX6850,WX6861,WX6851,WX6857,
    WX6854,WX6855,WX6858,WX6859,WX6864,WX6875,WX6865,WX6871,WX6868,WX6869,
    WX6872,WX6873,WX6878,WX6889,WX6879,WX6885,WX6882,WX6883,WX6886,WX6887,
    WX6892,WX6903,WX6893,WX6899,WX6896,WX6897,WX6900,WX6901,WX6906,WX6917,
    WX6907,WX6913,WX6910,WX6911,WX6914,WX6915,WX6920,WX6931,WX6921,WX6927,
    WX6924,WX6925,WX6928,WX6929,WX6934,WX6945,WX6935,WX6941,WX6938,WX6939,
    WX6942,WX6943,WX7472,WX7471,WX7473,WX7479,WX7478,WX7480,WX7486,WX7485,
    WX7487,WX7493,WX7492,WX7494,WX7500,WX7499,WX7501,WX7507,WX7506,WX7508,
    WX7514,WX7513,WX7515,WX7521,WX7520,WX7522,WX7528,WX7527,WX7529,WX7535,
    WX7534,WX7536,WX7542,WX7541,WX7543,WX7549,WX7548,WX7550,WX7556,WX7555,
    WX7557,WX7563,WX7562,WX7564,WX7570,WX7569,WX7571,WX7577,WX7576,WX7578,
    WX7584,WX7583,WX7585,WX7591,WX7590,WX7592,WX7598,WX7597,WX7599,WX7605,
    WX7604,WX7606,WX7612,WX7611,WX7613,WX7619,WX7618,WX7620,WX7626,WX7625,
    WX7627,WX7633,WX7632,WX7634,WX7640,WX7639,WX7641,WX7647,WX7646,WX7648,
    WX7654,WX7653,WX7655,WX7661,WX7660,WX7662,WX7668,WX7667,WX7669,WX7675,
    WX7674,WX7676,WX7682,WX7681,WX7683,WX7689,WX7688,WX7690,WX7699,WX7727,
    WX7726,WX7725,WX7698,WX7724,WX7723,WX7722,WX7721,WX7720,WX7719,WX7697,
    WX7718,WX7717,WX7716,WX7715,WX7696,WX7714,WX7713,WX7712,WX7711,WX7710,
    WX7709,WX7708,WX7707,WX7706,WX7705,WX7704,WX7703,WX7702,WX7701,WX7700,
    WX7793,WX7804,WX7794,WX7800,WX7797,WX7798,WX7801,WX7802,WX7807,WX7818,
    WX7808,WX7814,WX7811,WX7812,WX7815,WX7816,WX7821,WX7832,WX7822,WX7828,
    WX7825,WX7826,WX7829,WX7830,WX7835,WX7846,WX7836,WX7842,WX7839,WX7840,
    WX7843,WX7844,WX7849,WX7860,WX7850,WX7856,WX7853,WX7854,WX7857,WX7858,
    WX7863,WX7874,WX7864,WX7870,WX7867,WX7868,WX7871,WX7872,WX7877,WX7888,
    WX7878,WX7884,WX7881,WX7882,WX7885,WX7886,WX7891,WX7902,WX7892,WX7898,
    WX7895,WX7896,WX7899,WX7900,WX7905,WX7916,WX7906,WX7912,WX7909,WX7910,
    WX7913,WX7914,WX7919,WX7930,WX7920,WX7926,WX7923,WX7924,WX7927,WX7928,
    WX7933,WX7944,WX7934,WX7940,WX7937,WX7938,WX7941,WX7942,WX7947,WX7958,
    WX7948,WX7954,WX7951,WX7952,WX7955,WX7956,WX7961,WX7972,WX7962,WX7968,
    WX7965,WX7966,WX7969,WX7970,WX7975,WX7986,WX7976,WX7982,WX7979,WX7980,
    WX7983,WX7984,WX7989,WX8000,WX7990,WX7996,WX7993,WX7994,WX7997,WX7998,
    WX8003,WX8014,WX8004,WX8010,WX8007,WX8008,WX8011,WX8012,WX8017,WX8028,
    WX8018,WX8024,WX8021,WX8022,WX8025,WX8026,WX8031,WX8042,WX8032,WX8038,
    WX8035,WX8036,WX8039,WX8040,WX8045,WX8056,WX8046,WX8052,WX8049,WX8050,
    WX8053,WX8054,WX8059,WX8070,WX8060,WX8066,WX8063,WX8064,WX8067,WX8068,
    WX8073,WX8084,WX8074,WX8080,WX8077,WX8078,WX8081,WX8082,WX8087,WX8098,
    WX8088,WX8094,WX8091,WX8092,WX8095,WX8096,WX8101,WX8112,WX8102,WX8108,
    WX8105,WX8106,WX8109,WX8110,WX8115,WX8126,WX8116,WX8122,WX8119,WX8120,
    WX8123,WX8124,WX8129,WX8140,WX8130,WX8136,WX8133,WX8134,WX8137,WX8138,
    WX8143,WX8154,WX8144,WX8150,WX8147,WX8148,WX8151,WX8152,WX8157,WX8168,
    WX8158,WX8164,WX8161,WX8162,WX8165,WX8166,WX8171,WX8182,WX8172,WX8178,
    WX8175,WX8176,WX8179,WX8180,WX8185,WX8196,WX8186,WX8192,WX8189,WX8190,
    WX8193,WX8194,WX8199,WX8210,WX8200,WX8206,WX8203,WX8204,WX8207,WX8208,
    WX8213,WX8224,WX8214,WX8220,WX8217,WX8218,WX8221,WX8222,WX8227,WX8238,
    WX8228,WX8234,WX8231,WX8232,WX8235,WX8236,WX8765,WX8764,WX8766,WX8772,
    WX8771,WX8773,WX8779,WX8778,WX8780,WX8786,WX8785,WX8787,WX8793,WX8792,
    WX8794,WX8800,WX8799,WX8801,WX8807,WX8806,WX8808,WX8814,WX8813,WX8815,
    WX8821,WX8820,WX8822,WX8828,WX8827,WX8829,WX8835,WX8834,WX8836,WX8842,
    WX8841,WX8843,WX8849,WX8848,WX8850,WX8856,WX8855,WX8857,WX8863,WX8862,
    WX8864,WX8870,WX8869,WX8871,WX8877,WX8876,WX8878,WX8884,WX8883,WX8885,
    WX8891,WX8890,WX8892,WX8898,WX8897,WX8899,WX8905,WX8904,WX8906,WX8912,
    WX8911,WX8913,WX8919,WX8918,WX8920,WX8926,WX8925,WX8927,WX8933,WX8932,
    WX8934,WX8940,WX8939,WX8941,WX8947,WX8946,WX8948,WX8954,WX8953,WX8955,
    WX8961,WX8960,WX8962,WX8968,WX8967,WX8969,WX8975,WX8974,WX8976,WX8982,
    WX8981,WX8983,WX8992,WX9020,WX9019,WX9018,WX8991,WX9017,WX9016,WX9015,
    WX9014,WX9013,WX9012,WX8990,WX9011,WX9010,WX9009,WX9008,WX8989,WX9007,
    WX9006,WX9005,WX9004,WX9003,WX9002,WX9001,WX9000,WX8999,WX8998,WX8997,
    WX8996,WX8995,WX8994,WX8993,WX9086,WX9097,WX9087,WX9093,WX9090,WX9091,
    WX9094,WX9095,WX9100,WX9111,WX9101,WX9107,WX9104,WX9105,WX9108,WX9109,
    WX9114,WX9125,WX9115,WX9121,WX9118,WX9119,WX9122,WX9123,WX9128,WX9139,
    WX9129,WX9135,WX9132,WX9133,WX9136,WX9137,WX9142,WX9153,WX9143,WX9149,
    WX9146,WX9147,WX9150,WX9151,WX9156,WX9167,WX9157,WX9163,WX9160,WX9161,
    WX9164,WX9165,WX9170,WX9181,WX9171,WX9177,WX9174,WX9175,WX9178,WX9179,
    WX9184,WX9195,WX9185,WX9191,WX9188,WX9189,WX9192,WX9193,WX9198,WX9209,
    WX9199,WX9205,WX9202,WX9203,WX9206,WX9207,WX9212,WX9223,WX9213,WX9219,
    WX9216,WX9217,WX9220,WX9221,WX9226,WX9237,WX9227,WX9233,WX9230,WX9231,
    WX9234,WX9235,WX9240,WX9251,WX9241,WX9247,WX9244,WX9245,WX9248,WX9249,
    WX9254,WX9265,WX9255,WX9261,WX9258,WX9259,WX9262,WX9263,WX9268,WX9279,
    WX9269,WX9275,WX9272,WX9273,WX9276,WX9277,WX9282,WX9293,WX9283,WX9289,
    WX9286,WX9287,WX9290,WX9291,WX9296,WX9307,WX9297,WX9303,WX9300,WX9301,
    WX9304,WX9305,WX9310,WX9321,WX9311,WX9317,WX9314,WX9315,WX9318,WX9319,
    WX9324,WX9335,WX9325,WX9331,WX9328,WX9329,WX9332,WX9333,WX9338,WX9349,
    WX9339,WX9345,WX9342,WX9343,WX9346,WX9347,WX9352,WX9363,WX9353,WX9359,
    WX9356,WX9357,WX9360,WX9361,WX9366,WX9377,WX9367,WX9373,WX9370,WX9371,
    WX9374,WX9375,WX9380,WX9391,WX9381,WX9387,WX9384,WX9385,WX9388,WX9389,
    WX9394,WX9405,WX9395,WX9401,WX9398,WX9399,WX9402,WX9403,WX9408,WX9419,
    WX9409,WX9415,WX9412,WX9413,WX9416,WX9417,WX9422,WX9433,WX9423,WX9429,
    WX9426,WX9427,WX9430,WX9431,WX9436,WX9447,WX9437,WX9443,WX9440,WX9441,
    WX9444,WX9445,WX9450,WX9461,WX9451,WX9457,WX9454,WX9455,WX9458,WX9459,
    WX9464,WX9475,WX9465,WX9471,WX9468,WX9469,WX9472,WX9473,WX9478,WX9489,
    WX9479,WX9485,WX9482,WX9483,WX9486,WX9487,WX9492,WX9503,WX9493,WX9499,
    WX9496,WX9497,WX9500,WX9501,WX9506,WX9517,WX9507,WX9513,WX9510,WX9511,
    WX9514,WX9515,WX9520,WX9531,WX9521,WX9527,WX9524,WX9525,WX9528,WX9529,
    WX10058,WX10057,WX10059,WX10065,WX10064,WX10066,WX10072,WX10071,WX10073,
    WX10079,WX10078,WX10080,WX10086,WX10085,WX10087,WX10093,WX10092,WX10094,
    WX10100,WX10099,WX10101,WX10107,WX10106,WX10108,WX10114,WX10113,WX10115,
    WX10121,WX10120,WX10122,WX10128,WX10127,WX10129,WX10135,WX10134,WX10136,
    WX10142,WX10141,WX10143,WX10149,WX10148,WX10150,WX10156,WX10155,WX10157,
    WX10163,WX10162,WX10164,WX10170,WX10169,WX10171,WX10177,WX10176,WX10178,
    WX10184,WX10183,WX10185,WX10191,WX10190,WX10192,WX10198,WX10197,WX10199,
    WX10205,WX10204,WX10206,WX10212,WX10211,WX10213,WX10219,WX10218,WX10220,
    WX10226,WX10225,WX10227,WX10233,WX10232,WX10234,WX10240,WX10239,WX10241,
    WX10247,WX10246,WX10248,WX10254,WX10253,WX10255,WX10261,WX10260,WX10262,
    WX10268,WX10267,WX10269,WX10275,WX10274,WX10276,WX10285,WX10313,WX10312,
    WX10311,WX10284,WX10310,WX10309,WX10308,WX10307,WX10306,WX10305,WX10283,
    WX10304,WX10303,WX10302,WX10301,WX10282,WX10300,WX10299,WX10298,WX10297,
    WX10296,WX10295,WX10294,WX10293,WX10292,WX10291,WX10290,WX10289,WX10288,
    WX10287,WX10286,WX10379,WX10390,WX10380,WX10386,WX10383,WX10384,WX10387,
    WX10388,WX10393,WX10404,WX10394,WX10400,WX10397,WX10398,WX10401,WX10402,
    WX10407,WX10418,WX10408,WX10414,WX10411,WX10412,WX10415,WX10416,WX10421,
    WX10432,WX10422,WX10428,WX10425,WX10426,WX10429,WX10430,WX10435,WX10446,
    WX10436,WX10442,WX10439,WX10440,WX10443,WX10444,WX10449,WX10460,WX10450,
    WX10456,WX10453,WX10454,WX10457,WX10458,WX10463,WX10474,WX10464,WX10470,
    WX10467,WX10468,WX10471,WX10472,WX10477,WX10488,WX10478,WX10484,WX10481,
    WX10482,WX10485,WX10486,WX10491,WX10502,WX10492,WX10498,WX10495,WX10496,
    WX10499,WX10500,WX10505,WX10516,WX10506,WX10512,WX10509,WX10510,WX10513,
    WX10514,WX10519,WX10530,WX10520,WX10526,WX10523,WX10524,WX10527,WX10528,
    WX10533,WX10544,WX10534,WX10540,WX10537,WX10538,WX10541,WX10542,WX10547,
    WX10558,WX10548,WX10554,WX10551,WX10552,WX10555,WX10556,WX10561,WX10572,
    WX10562,WX10568,WX10565,WX10566,WX10569,WX10570,WX10575,WX10586,WX10576,
    WX10582,WX10579,WX10580,WX10583,WX10584,WX10589,WX10600,WX10590,WX10596,
    WX10593,WX10594,WX10597,WX10598,WX10603,WX10614,WX10604,WX10610,WX10607,
    WX10608,WX10611,WX10612,WX10617,WX10628,WX10618,WX10624,WX10621,WX10622,
    WX10625,WX10626,WX10631,WX10642,WX10632,WX10638,WX10635,WX10636,WX10639,
    WX10640,WX10645,WX10656,WX10646,WX10652,WX10649,WX10650,WX10653,WX10654,
    WX10659,WX10670,WX10660,WX10666,WX10663,WX10664,WX10667,WX10668,WX10673,
    WX10684,WX10674,WX10680,WX10677,WX10678,WX10681,WX10682,WX10687,WX10698,
    WX10688,WX10694,WX10691,WX10692,WX10695,WX10696,WX10701,WX10712,WX10702,
    WX10708,WX10705,WX10706,WX10709,WX10710,WX10715,WX10726,WX10716,WX10722,
    WX10719,WX10720,WX10723,WX10724,WX10729,WX10740,WX10730,WX10736,WX10733,
    WX10734,WX10737,WX10738,WX10743,WX10754,WX10744,WX10750,WX10747,WX10748,
    WX10751,WX10752,WX10757,WX10768,WX10758,WX10764,WX10761,WX10762,WX10765,
    WX10766,WX10771,WX10782,WX10772,WX10778,WX10775,WX10776,WX10779,WX10780,
    WX10785,WX10796,WX10786,WX10792,WX10789,WX10790,WX10793,WX10794,WX10799,
    WX10810,WX10800,WX10806,WX10803,WX10804,WX10807,WX10808,WX10813,WX10824,
    WX10814,WX10820,WX10817,WX10818,WX10821,WX10822,WX11351,WX11350,WX11352,
    WX11358,WX11357,WX11359,WX11365,WX11364,WX11366,WX11372,WX11371,WX11373,
    WX11379,WX11378,WX11380,WX11386,WX11385,WX11387,WX11393,WX11392,WX11394,
    WX11400,WX11399,WX11401,WX11407,WX11406,WX11408,WX11414,WX11413,WX11415,
    WX11421,WX11420,WX11422,WX11428,WX11427,WX11429,WX11435,WX11434,WX11436,
    WX11442,WX11441,WX11443,WX11449,WX11448,WX11450,WX11456,WX11455,WX11457,
    WX11463,WX11462,WX11464,WX11470,WX11469,WX11471,WX11477,WX11476,WX11478,
    WX11484,WX11483,WX11485,WX11491,WX11490,WX11492,WX11498,WX11497,WX11499,
    WX11505,WX11504,WX11506,WX11512,WX11511,WX11513,WX11519,WX11518,WX11520,
    WX11526,WX11525,WX11527,WX11533,WX11532,WX11534,WX11540,WX11539,WX11541,
    WX11547,WX11546,WX11548,WX11554,WX11553,WX11555,WX11561,WX11560,WX11562,
    WX11568,WX11567,WX11569,WX11578,WX11606,WX11605,WX11604,WX11577,WX11603,
    WX11602,WX11601,WX11600,WX11599,WX11598,WX11576,WX11597,WX11596,WX11595,
    WX11594,WX11575,WX11593,WX11592,WX11591,WX11590,WX11589,WX11588,WX11587,
    WX11586,WX11585,WX11584,WX11583,WX11582,WX11581,WX11580,WX11579,II1988,
    II1989,II1990,II1987,II1995,II1996,II1997,II1986,II2003,II2004,II2005,
    II2002,II2010,II2011,II2012,II2019,II2020,II2021,II2018,II2026,II2027,
    II2028,II2017,II2034,II2035,II2036,II2033,II2041,II2042,II2043,II2050,
    II2051,II2052,II2049,II2057,II2058,II2059,II2048,II2065,II2066,II2067,
    II2064,II2072,II2073,II2074,II2081,II2082,II2083,II2080,II2088,II2089,
    II2090,II2079,II2096,II2097,II2098,II2095,II2103,II2104,II2105,II2112,
    II2113,II2114,II2111,II2119,II2120,II2121,II2110,II2127,II2128,II2129,
    II2126,II2134,II2135,II2136,II2143,II2144,II2145,II2142,II2150,II2151,
    II2152,II2141,II2158,II2159,II2160,II2157,II2165,II2166,II2167,II2174,
    II2175,II2176,II2173,II2181,II2182,II2183,II2172,II2189,II2190,II2191,
    II2188,II2196,II2197,II2198,II2205,II2206,II2207,II2204,II2212,II2213,
    II2214,II2203,II2220,II2221,II2222,II2219,II2227,II2228,II2229,II2236,
    II2237,II2238,II2235,II2243,II2244,II2245,II2234,II2251,II2252,II2253,
    II2250,II2258,II2259,II2260,II2267,II2268,II2269,II2266,II2274,II2275,
    II2276,II2265,II2282,II2283,II2284,II2281,II2289,II2290,II2291,II2298,
    II2299,II2300,II2297,II2305,II2306,II2307,II2296,II2313,II2314,II2315,
    II2312,II2320,II2321,II2322,II2329,II2330,II2331,II2328,II2336,II2337,
    II2338,II2327,II2344,II2345,II2346,II2343,II2351,II2352,II2353,II2360,
    II2361,II2362,II2359,II2367,II2368,II2369,II2358,II2375,II2376,II2377,
    II2374,II2382,II2383,II2384,II2391,II2392,II2393,II2390,II2398,II2399,
    II2400,II2389,II2406,II2407,II2408,II2405,II2413,II2414,II2415,II2422,
    II2423,II2424,II2421,II2429,II2430,II2431,II2420,II2437,II2438,II2439,
    II2436,II2444,II2445,II2446,II2453,II2454,II2455,II2452,II2460,II2461,
    II2462,II2451,II2468,II2469,II2470,II2467,II2475,II2476,II2477,II2484,
    II2485,II2486,II2483,II2491,II2492,II2493,II2482,II2499,II2500,II2501,
    II2498,II2506,II2507,II2508,II2515,II2516,II2517,II2514,II2522,II2523,
    II2524,II2513,II2530,II2531,II2532,II2529,II2537,II2538,II2539,II2546,
    II2547,II2548,II2545,II2553,II2554,II2555,II2544,II2561,II2562,II2563,
    II2560,II2568,II2569,II2570,II2577,II2578,II2579,II2576,II2584,II2585,
    II2586,II2575,II2592,II2593,II2594,II2591,II2599,II2600,II2601,II2608,
    II2609,II2610,II2607,II2615,II2616,II2617,II2606,II2623,II2624,II2625,
    II2622,II2630,II2631,II2632,II2639,II2640,II2641,II2638,II2646,II2647,
    II2648,II2637,II2654,II2655,II2656,II2653,II2661,II2662,II2663,II2670,
    II2671,II2672,II2669,II2677,II2678,II2679,II2668,II2685,II2686,II2687,
    II2684,II2692,II2693,II2694,II2701,II2702,II2703,II2700,II2708,II2709,
    II2710,II2699,II2716,II2717,II2718,II2715,II2723,II2724,II2725,II2732,
    II2733,II2734,II2731,II2739,II2740,II2741,II2730,II2747,II2748,II2749,
    II2746,II2754,II2755,II2756,II2763,II2764,II2765,II2762,II2770,II2771,
    II2772,II2761,II2778,II2779,II2780,II2777,II2785,II2786,II2787,II2794,
    II2795,II2796,II2793,II2801,II2802,II2803,II2792,II2809,II2810,II2811,
    II2808,II2816,II2817,II2818,II2825,II2826,II2827,II2824,II2832,II2833,
    II2834,II2823,II2840,II2841,II2842,II2839,II2847,II2848,II2849,II2856,
    II2857,II2858,II2855,II2863,II2864,II2865,II2854,II2871,II2872,II2873,
    II2870,II2878,II2879,II2880,II2887,II2888,II2889,II2886,II2894,II2895,
    II2896,II2885,II2902,II2903,II2904,II2901,II2909,II2910,II2911,II2918,
    II2919,II2920,II2917,II2925,II2926,II2927,II2916,II2933,II2934,II2935,
    II2932,II2940,II2941,II2942,II2949,II2950,II2951,II2948,II2956,II2957,
    II2958,II2947,II2964,II2965,II2966,II2963,II2971,II2972,II2973,II3052,
    II3053,II3054,II3065,II3066,II3067,II3078,II3079,II3080,II3091,II3092,
    II3093,II3104,II3105,II3106,II3117,II3118,II3119,II3130,II3131,II3132,
    II3143,II3144,II3145,II3156,II3157,II3158,II3169,II3170,II3171,II3182,
    II3183,II3184,II3195,II3196,II3197,II3208,II3209,II3210,II3221,II3222,
    II3223,II3234,II3235,II3236,II3247,II3248,II3249,II3260,II3261,II3262,
    II3273,II3274,II3275,II3286,II3287,II3288,II3299,II3300,II3301,II3312,
    II3313,II3314,II3325,II3326,II3327,II3338,II3339,II3340,II3351,II3352,
    II3353,II3364,II3365,II3366,II3377,II3378,II3379,II3390,II3391,II3392,
    II3403,II3404,II3405,II3416,II3417,II3418,II3429,II3430,II3431,II3442,
    II3443,II3444,II3455,II3456,II3457,II3470,II3471,II3472,II3469,II3477,
    II3478,II3479,II3485,II3486,II3487,II3484,II3492,II3493,II3494,II3500,
    II3501,II3502,II3499,II3507,II3508,II3509,II3514,II3515,II3516,II3521,
    II3522,II3523,II3528,II3529,II3530,II3535,II3536,II3537,II3542,II3543,
    II3544,II3549,II3550,II3551,II3556,II3557,II3558,II3563,II3564,II3565,
    II3570,II3571,II3572,II3577,II3578,II3579,II3584,II3585,II3586,II3591,
    II3592,II3593,II3598,II3599,II3600,II3605,II3606,II3607,II3612,II3613,
    II3614,II3619,II3620,II3621,II3626,II3627,II3628,II3633,II3634,II3635,
    II3640,II3641,II3642,II3647,II3648,II3649,II3654,II3655,II3656,II3661,
    II3662,II3663,II3668,II3669,II3670,II3675,II3676,II3677,II3682,II3683,
    II3684,II3689,II3690,II3691,II3696,II3697,II3698,II3703,II3704,II3705,
    II3710,II3711,II3712,II5993,II5994,II5995,II5992,II6000,II6001,II6002,
    II5991,II6008,II6009,II6010,II6007,II6015,II6016,II6017,II6024,II6025,
    II6026,II6023,II6031,II6032,II6033,II6022,II6039,II6040,II6041,II6038,
    II6046,II6047,II6048,II6055,II6056,II6057,II6054,II6062,II6063,II6064,
    II6053,II6070,II6071,II6072,II6069,II6077,II6078,II6079,II6086,II6087,
    II6088,II6085,II6093,II6094,II6095,II6084,II6101,II6102,II6103,II6100,
    II6108,II6109,II6110,II6117,II6118,II6119,II6116,II6124,II6125,II6126,
    II6115,II6132,II6133,II6134,II6131,II6139,II6140,II6141,II6148,II6149,
    II6150,II6147,II6155,II6156,II6157,II6146,II6163,II6164,II6165,II6162,
    II6170,II6171,II6172,II6179,II6180,II6181,II6178,II6186,II6187,II6188,
    II6177,II6194,II6195,II6196,II6193,II6201,II6202,II6203,II6210,II6211,
    II6212,II6209,II6217,II6218,II6219,II6208,II6225,II6226,II6227,II6224,
    II6232,II6233,II6234,II6241,II6242,II6243,II6240,II6248,II6249,II6250,
    II6239,II6256,II6257,II6258,II6255,II6263,II6264,II6265,II6272,II6273,
    II6274,II6271,II6279,II6280,II6281,II6270,II6287,II6288,II6289,II6286,
    II6294,II6295,II6296,II6303,II6304,II6305,II6302,II6310,II6311,II6312,
    II6301,II6318,II6319,II6320,II6317,II6325,II6326,II6327,II6334,II6335,
    II6336,II6333,II6341,II6342,II6343,II6332,II6349,II6350,II6351,II6348,
    II6356,II6357,II6358,II6365,II6366,II6367,II6364,II6372,II6373,II6374,
    II6363,II6380,II6381,II6382,II6379,II6387,II6388,II6389,II6396,II6397,
    II6398,II6395,II6403,II6404,II6405,II6394,II6411,II6412,II6413,II6410,
    II6418,II6419,II6420,II6427,II6428,II6429,II6426,II6434,II6435,II6436,
    II6425,II6442,II6443,II6444,II6441,II6449,II6450,II6451,II6458,II6459,
    II6460,II6457,II6465,II6466,II6467,II6456,II6473,II6474,II6475,II6472,
    II6480,II6481,II6482,II6489,II6490,II6491,II6488,II6496,II6497,II6498,
    II6487,II6504,II6505,II6506,II6503,II6511,II6512,II6513,II6520,II6521,
    II6522,II6519,II6527,II6528,II6529,II6518,II6535,II6536,II6537,II6534,
    II6542,II6543,II6544,II6551,II6552,II6553,II6550,II6558,II6559,II6560,
    II6549,II6566,II6567,II6568,II6565,II6573,II6574,II6575,II6582,II6583,
    II6584,II6581,II6589,II6590,II6591,II6580,II6597,II6598,II6599,II6596,
    II6604,II6605,II6606,II6613,II6614,II6615,II6612,II6620,II6621,II6622,
    II6611,II6628,II6629,II6630,II6627,II6635,II6636,II6637,II6644,II6645,
    II6646,II6643,II6651,II6652,II6653,II6642,II6659,II6660,II6661,II6658,
    II6666,II6667,II6668,II6675,II6676,II6677,II6674,II6682,II6683,II6684,
    II6673,II6690,II6691,II6692,II6689,II6697,II6698,II6699,II6706,II6707,
    II6708,II6705,II6713,II6714,II6715,II6704,II6721,II6722,II6723,II6720,
    II6728,II6729,II6730,II6737,II6738,II6739,II6736,II6744,II6745,II6746,
    II6735,II6752,II6753,II6754,II6751,II6759,II6760,II6761,II6768,II6769,
    II6770,II6767,II6775,II6776,II6777,II6766,II6783,II6784,II6785,II6782,
    II6790,II6791,II6792,II6799,II6800,II6801,II6798,II6806,II6807,II6808,
    II6797,II6814,II6815,II6816,II6813,II6821,II6822,II6823,II6830,II6831,
    II6832,II6829,II6837,II6838,II6839,II6828,II6845,II6846,II6847,II6844,
    II6852,II6853,II6854,II6861,II6862,II6863,II6860,II6868,II6869,II6870,
    II6859,II6876,II6877,II6878,II6875,II6883,II6884,II6885,II6892,II6893,
    II6894,II6891,II6899,II6900,II6901,II6890,II6907,II6908,II6909,II6906,
    II6914,II6915,II6916,II6923,II6924,II6925,II6922,II6930,II6931,II6932,
    II6921,II6938,II6939,II6940,II6937,II6945,II6946,II6947,II6954,II6955,
    II6956,II6953,II6961,II6962,II6963,II6952,II6969,II6970,II6971,II6968,
    II6976,II6977,II6978,II7057,II7058,II7059,II7070,II7071,II7072,II7083,
    II7084,II7085,II7096,II7097,II7098,II7109,II7110,II7111,II7122,II7123,
    II7124,II7135,II7136,II7137,II7148,II7149,II7150,II7161,II7162,II7163,
    II7174,II7175,II7176,II7187,II7188,II7189,II7200,II7201,II7202,II7213,
    II7214,II7215,II7226,II7227,II7228,II7239,II7240,II7241,II7252,II7253,
    II7254,II7265,II7266,II7267,II7278,II7279,II7280,II7291,II7292,II7293,
    II7304,II7305,II7306,II7317,II7318,II7319,II7330,II7331,II7332,II7343,
    II7344,II7345,II7356,II7357,II7358,II7369,II7370,II7371,II7382,II7383,
    II7384,II7395,II7396,II7397,II7408,II7409,II7410,II7421,II7422,II7423,
    II7434,II7435,II7436,II7447,II7448,II7449,II7460,II7461,II7462,II7475,
    II7476,II7477,II7474,II7482,II7483,II7484,II7490,II7491,II7492,II7489,
    II7497,II7498,II7499,II7505,II7506,II7507,II7504,II7512,II7513,II7514,
    II7519,II7520,II7521,II7526,II7527,II7528,II7533,II7534,II7535,II7540,
    II7541,II7542,II7547,II7548,II7549,II7554,II7555,II7556,II7561,II7562,
    II7563,II7568,II7569,II7570,II7575,II7576,II7577,II7582,II7583,II7584,
    II7589,II7590,II7591,II7596,II7597,II7598,II7603,II7604,II7605,II7610,
    II7611,II7612,II7617,II7618,II7619,II7624,II7625,II7626,II7631,II7632,
    II7633,II7638,II7639,II7640,II7645,II7646,II7647,II7652,II7653,II7654,
    II7659,II7660,II7661,II7666,II7667,II7668,II7673,II7674,II7675,II7680,
    II7681,II7682,II7687,II7688,II7689,II7694,II7695,II7696,II7701,II7702,
    II7703,II7708,II7709,II7710,II7715,II7716,II7717,II9998,II9999,II10000,
    II9997,II10005,II10006,II10007,II9996,II10013,II10014,II10015,II10012,
    II10020,II10021,II10022,II10029,II10030,II10031,II10028,II10036,II10037,
    II10038,II10027,II10044,II10045,II10046,II10043,II10051,II10052,II10053,
    II10060,II10061,II10062,II10059,II10067,II10068,II10069,II10058,II10075,
    II10076,II10077,II10074,II10082,II10083,II10084,II10091,II10092,II10093,
    II10090,II10098,II10099,II10100,II10089,II10106,II10107,II10108,II10105,
    II10113,II10114,II10115,II10122,II10123,II10124,II10121,II10129,II10130,
    II10131,II10120,II10137,II10138,II10139,II10136,II10144,II10145,II10146,
    II10153,II10154,II10155,II10152,II10160,II10161,II10162,II10151,II10168,
    II10169,II10170,II10167,II10175,II10176,II10177,II10184,II10185,II10186,
    II10183,II10191,II10192,II10193,II10182,II10199,II10200,II10201,II10198,
    II10206,II10207,II10208,II10215,II10216,II10217,II10214,II10222,II10223,
    II10224,II10213,II10230,II10231,II10232,II10229,II10237,II10238,II10239,
    II10246,II10247,II10248,II10245,II10253,II10254,II10255,II10244,II10261,
    II10262,II10263,II10260,II10268,II10269,II10270,II10277,II10278,II10279,
    II10276,II10284,II10285,II10286,II10275,II10292,II10293,II10294,II10291,
    II10299,II10300,II10301,II10308,II10309,II10310,II10307,II10315,II10316,
    II10317,II10306,II10323,II10324,II10325,II10322,II10330,II10331,II10332,
    II10339,II10340,II10341,II10338,II10346,II10347,II10348,II10337,II10354,
    II10355,II10356,II10353,II10361,II10362,II10363,II10370,II10371,II10372,
    II10369,II10377,II10378,II10379,II10368,II10385,II10386,II10387,II10384,
    II10392,II10393,II10394,II10401,II10402,II10403,II10400,II10408,II10409,
    II10410,II10399,II10416,II10417,II10418,II10415,II10423,II10424,II10425,
    II10432,II10433,II10434,II10431,II10439,II10440,II10441,II10430,II10447,
    II10448,II10449,II10446,II10454,II10455,II10456,II10463,II10464,II10465,
    II10462,II10470,II10471,II10472,II10461,II10478,II10479,II10480,II10477,
    II10485,II10486,II10487,II10494,II10495,II10496,II10493,II10501,II10502,
    II10503,II10492,II10509,II10510,II10511,II10508,II10516,II10517,II10518,
    II10525,II10526,II10527,II10524,II10532,II10533,II10534,II10523,II10540,
    II10541,II10542,II10539,II10547,II10548,II10549,II10556,II10557,II10558,
    II10555,II10563,II10564,II10565,II10554,II10571,II10572,II10573,II10570,
    II10578,II10579,II10580,II10587,II10588,II10589,II10586,II10594,II10595,
    II10596,II10585,II10602,II10603,II10604,II10601,II10609,II10610,II10611,
    II10618,II10619,II10620,II10617,II10625,II10626,II10627,II10616,II10633,
    II10634,II10635,II10632,II10640,II10641,II10642,II10649,II10650,II10651,
    II10648,II10656,II10657,II10658,II10647,II10664,II10665,II10666,II10663,
    II10671,II10672,II10673,II10680,II10681,II10682,II10679,II10687,II10688,
    II10689,II10678,II10695,II10696,II10697,II10694,II10702,II10703,II10704,
    II10711,II10712,II10713,II10710,II10718,II10719,II10720,II10709,II10726,
    II10727,II10728,II10725,II10733,II10734,II10735,II10742,II10743,II10744,
    II10741,II10749,II10750,II10751,II10740,II10757,II10758,II10759,II10756,
    II10764,II10765,II10766,II10773,II10774,II10775,II10772,II10780,II10781,
    II10782,II10771,II10788,II10789,II10790,II10787,II10795,II10796,II10797,
    II10804,II10805,II10806,II10803,II10811,II10812,II10813,II10802,II10819,
    II10820,II10821,II10818,II10826,II10827,II10828,II10835,II10836,II10837,
    II10834,II10842,II10843,II10844,II10833,II10850,II10851,II10852,II10849,
    II10857,II10858,II10859,II10866,II10867,II10868,II10865,II10873,II10874,
    II10875,II10864,II10881,II10882,II10883,II10880,II10888,II10889,II10890,
    II10897,II10898,II10899,II10896,II10904,II10905,II10906,II10895,II10912,
    II10913,II10914,II10911,II10919,II10920,II10921,II10928,II10929,II10930,
    II10927,II10935,II10936,II10937,II10926,II10943,II10944,II10945,II10942,
    II10950,II10951,II10952,II10959,II10960,II10961,II10958,II10966,II10967,
    II10968,II10957,II10974,II10975,II10976,II10973,II10981,II10982,II10983,
    II11062,II11063,II11064,II11075,II11076,II11077,II11088,II11089,II11090,
    II11101,II11102,II11103,II11114,II11115,II11116,II11127,II11128,II11129,
    II11140,II11141,II11142,II11153,II11154,II11155,II11166,II11167,II11168,
    II11179,II11180,II11181,II11192,II11193,II11194,II11205,II11206,II11207,
    II11218,II11219,II11220,II11231,II11232,II11233,II11244,II11245,II11246,
    II11257,II11258,II11259,II11270,II11271,II11272,II11283,II11284,II11285,
    II11296,II11297,II11298,II11309,II11310,II11311,II11322,II11323,II11324,
    II11335,II11336,II11337,II11348,II11349,II11350,II11361,II11362,II11363,
    II11374,II11375,II11376,II11387,II11388,II11389,II11400,II11401,II11402,
    II11413,II11414,II11415,II11426,II11427,II11428,II11439,II11440,II11441,
    II11452,II11453,II11454,II11465,II11466,II11467,II11480,II11481,II11482,
    II11479,II11487,II11488,II11489,II11495,II11496,II11497,II11494,II11502,
    II11503,II11504,II11510,II11511,II11512,II11509,II11517,II11518,II11519,
    II11524,II11525,II11526,II11531,II11532,II11533,II11538,II11539,II11540,
    II11545,II11546,II11547,II11552,II11553,II11554,II11559,II11560,II11561,
    II11566,II11567,II11568,II11573,II11574,II11575,II11580,II11581,II11582,
    II11587,II11588,II11589,II11594,II11595,II11596,II11601,II11602,II11603,
    II11608,II11609,II11610,II11615,II11616,II11617,II11622,II11623,II11624,
    II11629,II11630,II11631,II11636,II11637,II11638,II11643,II11644,II11645,
    II11650,II11651,II11652,II11657,II11658,II11659,II11664,II11665,II11666,
    II11671,II11672,II11673,II11678,II11679,II11680,II11685,II11686,II11687,
    II11692,II11693,II11694,II11699,II11700,II11701,II11706,II11707,II11708,
    II11713,II11714,II11715,II11720,II11721,II11722,II14003,II14004,II14005,
    II14002,II14010,II14011,II14012,II14001,II14018,II14019,II14020,II14017,
    II14025,II14026,II14027,II14034,II14035,II14036,II14033,II14041,II14042,
    II14043,II14032,II14049,II14050,II14051,II14048,II14056,II14057,II14058,
    II14065,II14066,II14067,II14064,II14072,II14073,II14074,II14063,II14080,
    II14081,II14082,II14079,II14087,II14088,II14089,II14096,II14097,II14098,
    II14095,II14103,II14104,II14105,II14094,II14111,II14112,II14113,II14110,
    II14118,II14119,II14120,II14127,II14128,II14129,II14126,II14134,II14135,
    II14136,II14125,II14142,II14143,II14144,II14141,II14149,II14150,II14151,
    II14158,II14159,II14160,II14157,II14165,II14166,II14167,II14156,II14173,
    II14174,II14175,II14172,II14180,II14181,II14182,II14189,II14190,II14191,
    II14188,II14196,II14197,II14198,II14187,II14204,II14205,II14206,II14203,
    II14211,II14212,II14213,II14220,II14221,II14222,II14219,II14227,II14228,
    II14229,II14218,II14235,II14236,II14237,II14234,II14242,II14243,II14244,
    II14251,II14252,II14253,II14250,II14258,II14259,II14260,II14249,II14266,
    II14267,II14268,II14265,II14273,II14274,II14275,II14282,II14283,II14284,
    II14281,II14289,II14290,II14291,II14280,II14297,II14298,II14299,II14296,
    II14304,II14305,II14306,II14313,II14314,II14315,II14312,II14320,II14321,
    II14322,II14311,II14328,II14329,II14330,II14327,II14335,II14336,II14337,
    II14344,II14345,II14346,II14343,II14351,II14352,II14353,II14342,II14359,
    II14360,II14361,II14358,II14366,II14367,II14368,II14375,II14376,II14377,
    II14374,II14382,II14383,II14384,II14373,II14390,II14391,II14392,II14389,
    II14397,II14398,II14399,II14406,II14407,II14408,II14405,II14413,II14414,
    II14415,II14404,II14421,II14422,II14423,II14420,II14428,II14429,II14430,
    II14437,II14438,II14439,II14436,II14444,II14445,II14446,II14435,II14452,
    II14453,II14454,II14451,II14459,II14460,II14461,II14468,II14469,II14470,
    II14467,II14475,II14476,II14477,II14466,II14483,II14484,II14485,II14482,
    II14490,II14491,II14492,II14499,II14500,II14501,II14498,II14506,II14507,
    II14508,II14497,II14514,II14515,II14516,II14513,II14521,II14522,II14523,
    II14530,II14531,II14532,II14529,II14537,II14538,II14539,II14528,II14545,
    II14546,II14547,II14544,II14552,II14553,II14554,II14561,II14562,II14563,
    II14560,II14568,II14569,II14570,II14559,II14576,II14577,II14578,II14575,
    II14583,II14584,II14585,II14592,II14593,II14594,II14591,II14599,II14600,
    II14601,II14590,II14607,II14608,II14609,II14606,II14614,II14615,II14616,
    II14623,II14624,II14625,II14622,II14630,II14631,II14632,II14621,II14638,
    II14639,II14640,II14637,II14645,II14646,II14647,II14654,II14655,II14656,
    II14653,II14661,II14662,II14663,II14652,II14669,II14670,II14671,II14668,
    II14676,II14677,II14678,II14685,II14686,II14687,II14684,II14692,II14693,
    II14694,II14683,II14700,II14701,II14702,II14699,II14707,II14708,II14709,
    II14716,II14717,II14718,II14715,II14723,II14724,II14725,II14714,II14731,
    II14732,II14733,II14730,II14738,II14739,II14740,II14747,II14748,II14749,
    II14746,II14754,II14755,II14756,II14745,II14762,II14763,II14764,II14761,
    II14769,II14770,II14771,II14778,II14779,II14780,II14777,II14785,II14786,
    II14787,II14776,II14793,II14794,II14795,II14792,II14800,II14801,II14802,
    II14809,II14810,II14811,II14808,II14816,II14817,II14818,II14807,II14824,
    II14825,II14826,II14823,II14831,II14832,II14833,II14840,II14841,II14842,
    II14839,II14847,II14848,II14849,II14838,II14855,II14856,II14857,II14854,
    II14862,II14863,II14864,II14871,II14872,II14873,II14870,II14878,II14879,
    II14880,II14869,II14886,II14887,II14888,II14885,II14893,II14894,II14895,
    II14902,II14903,II14904,II14901,II14909,II14910,II14911,II14900,II14917,
    II14918,II14919,II14916,II14924,II14925,II14926,II14933,II14934,II14935,
    II14932,II14940,II14941,II14942,II14931,II14948,II14949,II14950,II14947,
    II14955,II14956,II14957,II14964,II14965,II14966,II14963,II14971,II14972,
    II14973,II14962,II14979,II14980,II14981,II14978,II14986,II14987,II14988,
    II15067,II15068,II15069,II15080,II15081,II15082,II15093,II15094,II15095,
    II15106,II15107,II15108,II15119,II15120,II15121,II15132,II15133,II15134,
    II15145,II15146,II15147,II15158,II15159,II15160,II15171,II15172,II15173,
    II15184,II15185,II15186,II15197,II15198,II15199,II15210,II15211,II15212,
    II15223,II15224,II15225,II15236,II15237,II15238,II15249,II15250,II15251,
    II15262,II15263,II15264,II15275,II15276,II15277,II15288,II15289,II15290,
    II15301,II15302,II15303,II15314,II15315,II15316,II15327,II15328,II15329,
    II15340,II15341,II15342,II15353,II15354,II15355,II15366,II15367,II15368,
    II15379,II15380,II15381,II15392,II15393,II15394,II15405,II15406,II15407,
    II15418,II15419,II15420,II15431,II15432,II15433,II15444,II15445,II15446,
    II15457,II15458,II15459,II15470,II15471,II15472,II15485,II15486,II15487,
    II15484,II15492,II15493,II15494,II15500,II15501,II15502,II15499,II15507,
    II15508,II15509,II15515,II15516,II15517,II15514,II15522,II15523,II15524,
    II15529,II15530,II15531,II15536,II15537,II15538,II15543,II15544,II15545,
    II15550,II15551,II15552,II15557,II15558,II15559,II15564,II15565,II15566,
    II15571,II15572,II15573,II15578,II15579,II15580,II15585,II15586,II15587,
    II15592,II15593,II15594,II15599,II15600,II15601,II15606,II15607,II15608,
    II15613,II15614,II15615,II15620,II15621,II15622,II15627,II15628,II15629,
    II15634,II15635,II15636,II15641,II15642,II15643,II15648,II15649,II15650,
    II15655,II15656,II15657,II15662,II15663,II15664,II15669,II15670,II15671,
    II15676,II15677,II15678,II15683,II15684,II15685,II15690,II15691,II15692,
    II15697,II15698,II15699,II15704,II15705,II15706,II15711,II15712,II15713,
    II15718,II15719,II15720,II15725,II15726,II15727,II18008,II18009,II18010,
    II18007,II18015,II18016,II18017,II18006,II18023,II18024,II18025,II18022,
    II18030,II18031,II18032,II18039,II18040,II18041,II18038,II18046,II18047,
    II18048,II18037,II18054,II18055,II18056,II18053,II18061,II18062,II18063,
    II18070,II18071,II18072,II18069,II18077,II18078,II18079,II18068,II18085,
    II18086,II18087,II18084,II18092,II18093,II18094,II18101,II18102,II18103,
    II18100,II18108,II18109,II18110,II18099,II18116,II18117,II18118,II18115,
    II18123,II18124,II18125,II18132,II18133,II18134,II18131,II18139,II18140,
    II18141,II18130,II18147,II18148,II18149,II18146,II18154,II18155,II18156,
    II18163,II18164,II18165,II18162,II18170,II18171,II18172,II18161,II18178,
    II18179,II18180,II18177,II18185,II18186,II18187,II18194,II18195,II18196,
    II18193,II18201,II18202,II18203,II18192,II18209,II18210,II18211,II18208,
    II18216,II18217,II18218,II18225,II18226,II18227,II18224,II18232,II18233,
    II18234,II18223,II18240,II18241,II18242,II18239,II18247,II18248,II18249,
    II18256,II18257,II18258,II18255,II18263,II18264,II18265,II18254,II18271,
    II18272,II18273,II18270,II18278,II18279,II18280,II18287,II18288,II18289,
    II18286,II18294,II18295,II18296,II18285,II18302,II18303,II18304,II18301,
    II18309,II18310,II18311,II18318,II18319,II18320,II18317,II18325,II18326,
    II18327,II18316,II18333,II18334,II18335,II18332,II18340,II18341,II18342,
    II18349,II18350,II18351,II18348,II18356,II18357,II18358,II18347,II18364,
    II18365,II18366,II18363,II18371,II18372,II18373,II18380,II18381,II18382,
    II18379,II18387,II18388,II18389,II18378,II18395,II18396,II18397,II18394,
    II18402,II18403,II18404,II18411,II18412,II18413,II18410,II18418,II18419,
    II18420,II18409,II18426,II18427,II18428,II18425,II18433,II18434,II18435,
    II18442,II18443,II18444,II18441,II18449,II18450,II18451,II18440,II18457,
    II18458,II18459,II18456,II18464,II18465,II18466,II18473,II18474,II18475,
    II18472,II18480,II18481,II18482,II18471,II18488,II18489,II18490,II18487,
    II18495,II18496,II18497,II18504,II18505,II18506,II18503,II18511,II18512,
    II18513,II18502,II18519,II18520,II18521,II18518,II18526,II18527,II18528,
    II18535,II18536,II18537,II18534,II18542,II18543,II18544,II18533,II18550,
    II18551,II18552,II18549,II18557,II18558,II18559,II18566,II18567,II18568,
    II18565,II18573,II18574,II18575,II18564,II18581,II18582,II18583,II18580,
    II18588,II18589,II18590,II18597,II18598,II18599,II18596,II18604,II18605,
    II18606,II18595,II18612,II18613,II18614,II18611,II18619,II18620,II18621,
    II18628,II18629,II18630,II18627,II18635,II18636,II18637,II18626,II18643,
    II18644,II18645,II18642,II18650,II18651,II18652,II18659,II18660,II18661,
    II18658,II18666,II18667,II18668,II18657,II18674,II18675,II18676,II18673,
    II18681,II18682,II18683,II18690,II18691,II18692,II18689,II18697,II18698,
    II18699,II18688,II18705,II18706,II18707,II18704,II18712,II18713,II18714,
    II18721,II18722,II18723,II18720,II18728,II18729,II18730,II18719,II18736,
    II18737,II18738,II18735,II18743,II18744,II18745,II18752,II18753,II18754,
    II18751,II18759,II18760,II18761,II18750,II18767,II18768,II18769,II18766,
    II18774,II18775,II18776,II18783,II18784,II18785,II18782,II18790,II18791,
    II18792,II18781,II18798,II18799,II18800,II18797,II18805,II18806,II18807,
    II18814,II18815,II18816,II18813,II18821,II18822,II18823,II18812,II18829,
    II18830,II18831,II18828,II18836,II18837,II18838,II18845,II18846,II18847,
    II18844,II18852,II18853,II18854,II18843,II18860,II18861,II18862,II18859,
    II18867,II18868,II18869,II18876,II18877,II18878,II18875,II18883,II18884,
    II18885,II18874,II18891,II18892,II18893,II18890,II18898,II18899,II18900,
    II18907,II18908,II18909,II18906,II18914,II18915,II18916,II18905,II18922,
    II18923,II18924,II18921,II18929,II18930,II18931,II18938,II18939,II18940,
    II18937,II18945,II18946,II18947,II18936,II18953,II18954,II18955,II18952,
    II18960,II18961,II18962,II18969,II18970,II18971,II18968,II18976,II18977,
    II18978,II18967,II18984,II18985,II18986,II18983,II18991,II18992,II18993,
    II19072,II19073,II19074,II19085,II19086,II19087,II19098,II19099,II19100,
    II19111,II19112,II19113,II19124,II19125,II19126,II19137,II19138,II19139,
    II19150,II19151,II19152,II19163,II19164,II19165,II19176,II19177,II19178,
    II19189,II19190,II19191,II19202,II19203,II19204,II19215,II19216,II19217,
    II19228,II19229,II19230,II19241,II19242,II19243,II19254,II19255,II19256,
    II19267,II19268,II19269,II19280,II19281,II19282,II19293,II19294,II19295,
    II19306,II19307,II19308,II19319,II19320,II19321,II19332,II19333,II19334,
    II19345,II19346,II19347,II19358,II19359,II19360,II19371,II19372,II19373,
    II19384,II19385,II19386,II19397,II19398,II19399,II19410,II19411,II19412,
    II19423,II19424,II19425,II19436,II19437,II19438,II19449,II19450,II19451,
    II19462,II19463,II19464,II19475,II19476,II19477,II19490,II19491,II19492,
    II19489,II19497,II19498,II19499,II19505,II19506,II19507,II19504,II19512,
    II19513,II19514,II19520,II19521,II19522,II19519,II19527,II19528,II19529,
    II19534,II19535,II19536,II19541,II19542,II19543,II19548,II19549,II19550,
    II19555,II19556,II19557,II19562,II19563,II19564,II19569,II19570,II19571,
    II19576,II19577,II19578,II19583,II19584,II19585,II19590,II19591,II19592,
    II19597,II19598,II19599,II19604,II19605,II19606,II19611,II19612,II19613,
    II19618,II19619,II19620,II19625,II19626,II19627,II19632,II19633,II19634,
    II19639,II19640,II19641,II19646,II19647,II19648,II19653,II19654,II19655,
    II19660,II19661,II19662,II19667,II19668,II19669,II19674,II19675,II19676,
    II19681,II19682,II19683,II19688,II19689,II19690,II19695,II19696,II19697,
    II19702,II19703,II19704,II19709,II19710,II19711,II19716,II19717,II19718,
    II19723,II19724,II19725,II19730,II19731,II19732,II22013,II22014,II22015,
    II22012,II22020,II22021,II22022,II22011,II22028,II22029,II22030,II22027,
    II22035,II22036,II22037,II22044,II22045,II22046,II22043,II22051,II22052,
    II22053,II22042,II22059,II22060,II22061,II22058,II22066,II22067,II22068,
    II22075,II22076,II22077,II22074,II22082,II22083,II22084,II22073,II22090,
    II22091,II22092,II22089,II22097,II22098,II22099,II22106,II22107,II22108,
    II22105,II22113,II22114,II22115,II22104,II22121,II22122,II22123,II22120,
    II22128,II22129,II22130,II22137,II22138,II22139,II22136,II22144,II22145,
    II22146,II22135,II22152,II22153,II22154,II22151,II22159,II22160,II22161,
    II22168,II22169,II22170,II22167,II22175,II22176,II22177,II22166,II22183,
    II22184,II22185,II22182,II22190,II22191,II22192,II22199,II22200,II22201,
    II22198,II22206,II22207,II22208,II22197,II22214,II22215,II22216,II22213,
    II22221,II22222,II22223,II22230,II22231,II22232,II22229,II22237,II22238,
    II22239,II22228,II22245,II22246,II22247,II22244,II22252,II22253,II22254,
    II22261,II22262,II22263,II22260,II22268,II22269,II22270,II22259,II22276,
    II22277,II22278,II22275,II22283,II22284,II22285,II22292,II22293,II22294,
    II22291,II22299,II22300,II22301,II22290,II22307,II22308,II22309,II22306,
    II22314,II22315,II22316,II22323,II22324,II22325,II22322,II22330,II22331,
    II22332,II22321,II22338,II22339,II22340,II22337,II22345,II22346,II22347,
    II22354,II22355,II22356,II22353,II22361,II22362,II22363,II22352,II22369,
    II22370,II22371,II22368,II22376,II22377,II22378,II22385,II22386,II22387,
    II22384,II22392,II22393,II22394,II22383,II22400,II22401,II22402,II22399,
    II22407,II22408,II22409,II22416,II22417,II22418,II22415,II22423,II22424,
    II22425,II22414,II22431,II22432,II22433,II22430,II22438,II22439,II22440,
    II22447,II22448,II22449,II22446,II22454,II22455,II22456,II22445,II22462,
    II22463,II22464,II22461,II22469,II22470,II22471,II22478,II22479,II22480,
    II22477,II22485,II22486,II22487,II22476,II22493,II22494,II22495,II22492,
    II22500,II22501,II22502,II22509,II22510,II22511,II22508,II22516,II22517,
    II22518,II22507,II22524,II22525,II22526,II22523,II22531,II22532,II22533,
    II22540,II22541,II22542,II22539,II22547,II22548,II22549,II22538,II22555,
    II22556,II22557,II22554,II22562,II22563,II22564,II22571,II22572,II22573,
    II22570,II22578,II22579,II22580,II22569,II22586,II22587,II22588,II22585,
    II22593,II22594,II22595,II22602,II22603,II22604,II22601,II22609,II22610,
    II22611,II22600,II22617,II22618,II22619,II22616,II22624,II22625,II22626,
    II22633,II22634,II22635,II22632,II22640,II22641,II22642,II22631,II22648,
    II22649,II22650,II22647,II22655,II22656,II22657,II22664,II22665,II22666,
    II22663,II22671,II22672,II22673,II22662,II22679,II22680,II22681,II22678,
    II22686,II22687,II22688,II22695,II22696,II22697,II22694,II22702,II22703,
    II22704,II22693,II22710,II22711,II22712,II22709,II22717,II22718,II22719,
    II22726,II22727,II22728,II22725,II22733,II22734,II22735,II22724,II22741,
    II22742,II22743,II22740,II22748,II22749,II22750,II22757,II22758,II22759,
    II22756,II22764,II22765,II22766,II22755,II22772,II22773,II22774,II22771,
    II22779,II22780,II22781,II22788,II22789,II22790,II22787,II22795,II22796,
    II22797,II22786,II22803,II22804,II22805,II22802,II22810,II22811,II22812,
    II22819,II22820,II22821,II22818,II22826,II22827,II22828,II22817,II22834,
    II22835,II22836,II22833,II22841,II22842,II22843,II22850,II22851,II22852,
    II22849,II22857,II22858,II22859,II22848,II22865,II22866,II22867,II22864,
    II22872,II22873,II22874,II22881,II22882,II22883,II22880,II22888,II22889,
    II22890,II22879,II22896,II22897,II22898,II22895,II22903,II22904,II22905,
    II22912,II22913,II22914,II22911,II22919,II22920,II22921,II22910,II22927,
    II22928,II22929,II22926,II22934,II22935,II22936,II22943,II22944,II22945,
    II22942,II22950,II22951,II22952,II22941,II22958,II22959,II22960,II22957,
    II22965,II22966,II22967,II22974,II22975,II22976,II22973,II22981,II22982,
    II22983,II22972,II22989,II22990,II22991,II22988,II22996,II22997,II22998,
    II23077,II23078,II23079,II23090,II23091,II23092,II23103,II23104,II23105,
    II23116,II23117,II23118,II23129,II23130,II23131,II23142,II23143,II23144,
    II23155,II23156,II23157,II23168,II23169,II23170,II23181,II23182,II23183,
    II23194,II23195,II23196,II23207,II23208,II23209,II23220,II23221,II23222,
    II23233,II23234,II23235,II23246,II23247,II23248,II23259,II23260,II23261,
    II23272,II23273,II23274,II23285,II23286,II23287,II23298,II23299,II23300,
    II23311,II23312,II23313,II23324,II23325,II23326,II23337,II23338,II23339,
    II23350,II23351,II23352,II23363,II23364,II23365,II23376,II23377,II23378,
    II23389,II23390,II23391,II23402,II23403,II23404,II23415,II23416,II23417,
    II23428,II23429,II23430,II23441,II23442,II23443,II23454,II23455,II23456,
    II23467,II23468,II23469,II23480,II23481,II23482,II23495,II23496,II23497,
    II23494,II23502,II23503,II23504,II23510,II23511,II23512,II23509,II23517,
    II23518,II23519,II23525,II23526,II23527,II23524,II23532,II23533,II23534,
    II23539,II23540,II23541,II23546,II23547,II23548,II23553,II23554,II23555,
    II23560,II23561,II23562,II23567,II23568,II23569,II23574,II23575,II23576,
    II23581,II23582,II23583,II23588,II23589,II23590,II23595,II23596,II23597,
    II23602,II23603,II23604,II23609,II23610,II23611,II23616,II23617,II23618,
    II23623,II23624,II23625,II23630,II23631,II23632,II23637,II23638,II23639,
    II23644,II23645,II23646,II23651,II23652,II23653,II23658,II23659,II23660,
    II23665,II23666,II23667,II23672,II23673,II23674,II23679,II23680,II23681,
    II23686,II23687,II23688,II23693,II23694,II23695,II23700,II23701,II23702,
    II23707,II23708,II23709,II23714,II23715,II23716,II23721,II23722,II23723,
    II23728,II23729,II23730,II23735,II23736,II23737,II26018,II26019,II26020,
    II26017,II26025,II26026,II26027,II26016,II26033,II26034,II26035,II26032,
    II26040,II26041,II26042,II26049,II26050,II26051,II26048,II26056,II26057,
    II26058,II26047,II26064,II26065,II26066,II26063,II26071,II26072,II26073,
    II26080,II26081,II26082,II26079,II26087,II26088,II26089,II26078,II26095,
    II26096,II26097,II26094,II26102,II26103,II26104,II26111,II26112,II26113,
    II26110,II26118,II26119,II26120,II26109,II26126,II26127,II26128,II26125,
    II26133,II26134,II26135,II26142,II26143,II26144,II26141,II26149,II26150,
    II26151,II26140,II26157,II26158,II26159,II26156,II26164,II26165,II26166,
    II26173,II26174,II26175,II26172,II26180,II26181,II26182,II26171,II26188,
    II26189,II26190,II26187,II26195,II26196,II26197,II26204,II26205,II26206,
    II26203,II26211,II26212,II26213,II26202,II26219,II26220,II26221,II26218,
    II26226,II26227,II26228,II26235,II26236,II26237,II26234,II26242,II26243,
    II26244,II26233,II26250,II26251,II26252,II26249,II26257,II26258,II26259,
    II26266,II26267,II26268,II26265,II26273,II26274,II26275,II26264,II26281,
    II26282,II26283,II26280,II26288,II26289,II26290,II26297,II26298,II26299,
    II26296,II26304,II26305,II26306,II26295,II26312,II26313,II26314,II26311,
    II26319,II26320,II26321,II26328,II26329,II26330,II26327,II26335,II26336,
    II26337,II26326,II26343,II26344,II26345,II26342,II26350,II26351,II26352,
    II26359,II26360,II26361,II26358,II26366,II26367,II26368,II26357,II26374,
    II26375,II26376,II26373,II26381,II26382,II26383,II26390,II26391,II26392,
    II26389,II26397,II26398,II26399,II26388,II26405,II26406,II26407,II26404,
    II26412,II26413,II26414,II26421,II26422,II26423,II26420,II26428,II26429,
    II26430,II26419,II26436,II26437,II26438,II26435,II26443,II26444,II26445,
    II26452,II26453,II26454,II26451,II26459,II26460,II26461,II26450,II26467,
    II26468,II26469,II26466,II26474,II26475,II26476,II26483,II26484,II26485,
    II26482,II26490,II26491,II26492,II26481,II26498,II26499,II26500,II26497,
    II26505,II26506,II26507,II26514,II26515,II26516,II26513,II26521,II26522,
    II26523,II26512,II26529,II26530,II26531,II26528,II26536,II26537,II26538,
    II26545,II26546,II26547,II26544,II26552,II26553,II26554,II26543,II26560,
    II26561,II26562,II26559,II26567,II26568,II26569,II26576,II26577,II26578,
    II26575,II26583,II26584,II26585,II26574,II26591,II26592,II26593,II26590,
    II26598,II26599,II26600,II26607,II26608,II26609,II26606,II26614,II26615,
    II26616,II26605,II26622,II26623,II26624,II26621,II26629,II26630,II26631,
    II26638,II26639,II26640,II26637,II26645,II26646,II26647,II26636,II26653,
    II26654,II26655,II26652,II26660,II26661,II26662,II26669,II26670,II26671,
    II26668,II26676,II26677,II26678,II26667,II26684,II26685,II26686,II26683,
    II26691,II26692,II26693,II26700,II26701,II26702,II26699,II26707,II26708,
    II26709,II26698,II26715,II26716,II26717,II26714,II26722,II26723,II26724,
    II26731,II26732,II26733,II26730,II26738,II26739,II26740,II26729,II26746,
    II26747,II26748,II26745,II26753,II26754,II26755,II26762,II26763,II26764,
    II26761,II26769,II26770,II26771,II26760,II26777,II26778,II26779,II26776,
    II26784,II26785,II26786,II26793,II26794,II26795,II26792,II26800,II26801,
    II26802,II26791,II26808,II26809,II26810,II26807,II26815,II26816,II26817,
    II26824,II26825,II26826,II26823,II26831,II26832,II26833,II26822,II26839,
    II26840,II26841,II26838,II26846,II26847,II26848,II26855,II26856,II26857,
    II26854,II26862,II26863,II26864,II26853,II26870,II26871,II26872,II26869,
    II26877,II26878,II26879,II26886,II26887,II26888,II26885,II26893,II26894,
    II26895,II26884,II26901,II26902,II26903,II26900,II26908,II26909,II26910,
    II26917,II26918,II26919,II26916,II26924,II26925,II26926,II26915,II26932,
    II26933,II26934,II26931,II26939,II26940,II26941,II26948,II26949,II26950,
    II26947,II26955,II26956,II26957,II26946,II26963,II26964,II26965,II26962,
    II26970,II26971,II26972,II26979,II26980,II26981,II26978,II26986,II26987,
    II26988,II26977,II26994,II26995,II26996,II26993,II27001,II27002,II27003,
    II27082,II27083,II27084,II27095,II27096,II27097,II27108,II27109,II27110,
    II27121,II27122,II27123,II27134,II27135,II27136,II27147,II27148,II27149,
    II27160,II27161,II27162,II27173,II27174,II27175,II27186,II27187,II27188,
    II27199,II27200,II27201,II27212,II27213,II27214,II27225,II27226,II27227,
    II27238,II27239,II27240,II27251,II27252,II27253,II27264,II27265,II27266,
    II27277,II27278,II27279,II27290,II27291,II27292,II27303,II27304,II27305,
    II27316,II27317,II27318,II27329,II27330,II27331,II27342,II27343,II27344,
    II27355,II27356,II27357,II27368,II27369,II27370,II27381,II27382,II27383,
    II27394,II27395,II27396,II27407,II27408,II27409,II27420,II27421,II27422,
    II27433,II27434,II27435,II27446,II27447,II27448,II27459,II27460,II27461,
    II27472,II27473,II27474,II27485,II27486,II27487,II27500,II27501,II27502,
    II27499,II27507,II27508,II27509,II27515,II27516,II27517,II27514,II27522,
    II27523,II27524,II27530,II27531,II27532,II27529,II27537,II27538,II27539,
    II27544,II27545,II27546,II27551,II27552,II27553,II27558,II27559,II27560,
    II27565,II27566,II27567,II27572,II27573,II27574,II27579,II27580,II27581,
    II27586,II27587,II27588,II27593,II27594,II27595,II27600,II27601,II27602,
    II27607,II27608,II27609,II27614,II27615,II27616,II27621,II27622,II27623,
    II27628,II27629,II27630,II27635,II27636,II27637,II27642,II27643,II27644,
    II27649,II27650,II27651,II27656,II27657,II27658,II27663,II27664,II27665,
    II27670,II27671,II27672,II27677,II27678,II27679,II27684,II27685,II27686,
    II27691,II27692,II27693,II27698,II27699,II27700,II27705,II27706,II27707,
    II27712,II27713,II27714,II27719,II27720,II27721,II27726,II27727,II27728,
    II27733,II27734,II27735,II27740,II27741,II27742,II30023,II30024,II30025,
    II30022,II30030,II30031,II30032,II30021,II30038,II30039,II30040,II30037,
    II30045,II30046,II30047,II30054,II30055,II30056,II30053,II30061,II30062,
    II30063,II30052,II30069,II30070,II30071,II30068,II30076,II30077,II30078,
    II30085,II30086,II30087,II30084,II30092,II30093,II30094,II30083,II30100,
    II30101,II30102,II30099,II30107,II30108,II30109,II30116,II30117,II30118,
    II30115,II30123,II30124,II30125,II30114,II30131,II30132,II30133,II30130,
    II30138,II30139,II30140,II30147,II30148,II30149,II30146,II30154,II30155,
    II30156,II30145,II30162,II30163,II30164,II30161,II30169,II30170,II30171,
    II30178,II30179,II30180,II30177,II30185,II30186,II30187,II30176,II30193,
    II30194,II30195,II30192,II30200,II30201,II30202,II30209,II30210,II30211,
    II30208,II30216,II30217,II30218,II30207,II30224,II30225,II30226,II30223,
    II30231,II30232,II30233,II30240,II30241,II30242,II30239,II30247,II30248,
    II30249,II30238,II30255,II30256,II30257,II30254,II30262,II30263,II30264,
    II30271,II30272,II30273,II30270,II30278,II30279,II30280,II30269,II30286,
    II30287,II30288,II30285,II30293,II30294,II30295,II30302,II30303,II30304,
    II30301,II30309,II30310,II30311,II30300,II30317,II30318,II30319,II30316,
    II30324,II30325,II30326,II30333,II30334,II30335,II30332,II30340,II30341,
    II30342,II30331,II30348,II30349,II30350,II30347,II30355,II30356,II30357,
    II30364,II30365,II30366,II30363,II30371,II30372,II30373,II30362,II30379,
    II30380,II30381,II30378,II30386,II30387,II30388,II30395,II30396,II30397,
    II30394,II30402,II30403,II30404,II30393,II30410,II30411,II30412,II30409,
    II30417,II30418,II30419,II30426,II30427,II30428,II30425,II30433,II30434,
    II30435,II30424,II30441,II30442,II30443,II30440,II30448,II30449,II30450,
    II30457,II30458,II30459,II30456,II30464,II30465,II30466,II30455,II30472,
    II30473,II30474,II30471,II30479,II30480,II30481,II30488,II30489,II30490,
    II30487,II30495,II30496,II30497,II30486,II30503,II30504,II30505,II30502,
    II30510,II30511,II30512,II30519,II30520,II30521,II30518,II30526,II30527,
    II30528,II30517,II30534,II30535,II30536,II30533,II30541,II30542,II30543,
    II30550,II30551,II30552,II30549,II30557,II30558,II30559,II30548,II30565,
    II30566,II30567,II30564,II30572,II30573,II30574,II30581,II30582,II30583,
    II30580,II30588,II30589,II30590,II30579,II30596,II30597,II30598,II30595,
    II30603,II30604,II30605,II30612,II30613,II30614,II30611,II30619,II30620,
    II30621,II30610,II30627,II30628,II30629,II30626,II30634,II30635,II30636,
    II30643,II30644,II30645,II30642,II30650,II30651,II30652,II30641,II30658,
    II30659,II30660,II30657,II30665,II30666,II30667,II30674,II30675,II30676,
    II30673,II30681,II30682,II30683,II30672,II30689,II30690,II30691,II30688,
    II30696,II30697,II30698,II30705,II30706,II30707,II30704,II30712,II30713,
    II30714,II30703,II30720,II30721,II30722,II30719,II30727,II30728,II30729,
    II30736,II30737,II30738,II30735,II30743,II30744,II30745,II30734,II30751,
    II30752,II30753,II30750,II30758,II30759,II30760,II30767,II30768,II30769,
    II30766,II30774,II30775,II30776,II30765,II30782,II30783,II30784,II30781,
    II30789,II30790,II30791,II30798,II30799,II30800,II30797,II30805,II30806,
    II30807,II30796,II30813,II30814,II30815,II30812,II30820,II30821,II30822,
    II30829,II30830,II30831,II30828,II30836,II30837,II30838,II30827,II30844,
    II30845,II30846,II30843,II30851,II30852,II30853,II30860,II30861,II30862,
    II30859,II30867,II30868,II30869,II30858,II30875,II30876,II30877,II30874,
    II30882,II30883,II30884,II30891,II30892,II30893,II30890,II30898,II30899,
    II30900,II30889,II30906,II30907,II30908,II30905,II30913,II30914,II30915,
    II30922,II30923,II30924,II30921,II30929,II30930,II30931,II30920,II30937,
    II30938,II30939,II30936,II30944,II30945,II30946,II30953,II30954,II30955,
    II30952,II30960,II30961,II30962,II30951,II30968,II30969,II30970,II30967,
    II30975,II30976,II30977,II30984,II30985,II30986,II30983,II30991,II30992,
    II30993,II30982,II30999,II31000,II31001,II30998,II31006,II31007,II31008,
    II31087,II31088,II31089,II31100,II31101,II31102,II31113,II31114,II31115,
    II31126,II31127,II31128,II31139,II31140,II31141,II31152,II31153,II31154,
    II31165,II31166,II31167,II31178,II31179,II31180,II31191,II31192,II31193,
    II31204,II31205,II31206,II31217,II31218,II31219,II31230,II31231,II31232,
    II31243,II31244,II31245,II31256,II31257,II31258,II31269,II31270,II31271,
    II31282,II31283,II31284,II31295,II31296,II31297,II31308,II31309,II31310,
    II31321,II31322,II31323,II31334,II31335,II31336,II31347,II31348,II31349,
    II31360,II31361,II31362,II31373,II31374,II31375,II31386,II31387,II31388,
    II31399,II31400,II31401,II31412,II31413,II31414,II31425,II31426,II31427,
    II31438,II31439,II31440,II31451,II31452,II31453,II31464,II31465,II31466,
    II31477,II31478,II31479,II31490,II31491,II31492,II31505,II31506,II31507,
    II31504,II31512,II31513,II31514,II31520,II31521,II31522,II31519,II31527,
    II31528,II31529,II31535,II31536,II31537,II31534,II31542,II31543,II31544,
    II31549,II31550,II31551,II31556,II31557,II31558,II31563,II31564,II31565,
    II31570,II31571,II31572,II31577,II31578,II31579,II31584,II31585,II31586,
    II31591,II31592,II31593,II31598,II31599,II31600,II31605,II31606,II31607,
    II31612,II31613,II31614,II31619,II31620,II31621,II31626,II31627,II31628,
    II31633,II31634,II31635,II31640,II31641,II31642,II31647,II31648,II31649,
    II31654,II31655,II31656,II31661,II31662,II31663,II31668,II31669,II31670,
    II31675,II31676,II31677,II31682,II31683,II31684,II31689,II31690,II31691,
    II31696,II31697,II31698,II31703,II31704,II31705,II31710,II31711,II31712,
    II31717,II31718,II31719,II31724,II31725,II31726,II31731,II31732,II31733,
    II31738,II31739,II31740,II31745,II31746,II31747,II34028,II34029,II34030,
    II34027,II34035,II34036,II34037,II34026,II34043,II34044,II34045,II34042,
    II34050,II34051,II34052,II34059,II34060,II34061,II34058,II34066,II34067,
    II34068,II34057,II34074,II34075,II34076,II34073,II34081,II34082,II34083,
    II34090,II34091,II34092,II34089,II34097,II34098,II34099,II34088,II34105,
    II34106,II34107,II34104,II34112,II34113,II34114,II34121,II34122,II34123,
    II34120,II34128,II34129,II34130,II34119,II34136,II34137,II34138,II34135,
    II34143,II34144,II34145,II34152,II34153,II34154,II34151,II34159,II34160,
    II34161,II34150,II34167,II34168,II34169,II34166,II34174,II34175,II34176,
    II34183,II34184,II34185,II34182,II34190,II34191,II34192,II34181,II34198,
    II34199,II34200,II34197,II34205,II34206,II34207,II34214,II34215,II34216,
    II34213,II34221,II34222,II34223,II34212,II34229,II34230,II34231,II34228,
    II34236,II34237,II34238,II34245,II34246,II34247,II34244,II34252,II34253,
    II34254,II34243,II34260,II34261,II34262,II34259,II34267,II34268,II34269,
    II34276,II34277,II34278,II34275,II34283,II34284,II34285,II34274,II34291,
    II34292,II34293,II34290,II34298,II34299,II34300,II34307,II34308,II34309,
    II34306,II34314,II34315,II34316,II34305,II34322,II34323,II34324,II34321,
    II34329,II34330,II34331,II34338,II34339,II34340,II34337,II34345,II34346,
    II34347,II34336,II34353,II34354,II34355,II34352,II34360,II34361,II34362,
    II34369,II34370,II34371,II34368,II34376,II34377,II34378,II34367,II34384,
    II34385,II34386,II34383,II34391,II34392,II34393,II34400,II34401,II34402,
    II34399,II34407,II34408,II34409,II34398,II34415,II34416,II34417,II34414,
    II34422,II34423,II34424,II34431,II34432,II34433,II34430,II34438,II34439,
    II34440,II34429,II34446,II34447,II34448,II34445,II34453,II34454,II34455,
    II34462,II34463,II34464,II34461,II34469,II34470,II34471,II34460,II34477,
    II34478,II34479,II34476,II34484,II34485,II34486,II34493,II34494,II34495,
    II34492,II34500,II34501,II34502,II34491,II34508,II34509,II34510,II34507,
    II34515,II34516,II34517,II34524,II34525,II34526,II34523,II34531,II34532,
    II34533,II34522,II34539,II34540,II34541,II34538,II34546,II34547,II34548,
    II34555,II34556,II34557,II34554,II34562,II34563,II34564,II34553,II34570,
    II34571,II34572,II34569,II34577,II34578,II34579,II34586,II34587,II34588,
    II34585,II34593,II34594,II34595,II34584,II34601,II34602,II34603,II34600,
    II34608,II34609,II34610,II34617,II34618,II34619,II34616,II34624,II34625,
    II34626,II34615,II34632,II34633,II34634,II34631,II34639,II34640,II34641,
    II34648,II34649,II34650,II34647,II34655,II34656,II34657,II34646,II34663,
    II34664,II34665,II34662,II34670,II34671,II34672,II34679,II34680,II34681,
    II34678,II34686,II34687,II34688,II34677,II34694,II34695,II34696,II34693,
    II34701,II34702,II34703,II34710,II34711,II34712,II34709,II34717,II34718,
    II34719,II34708,II34725,II34726,II34727,II34724,II34732,II34733,II34734,
    II34741,II34742,II34743,II34740,II34748,II34749,II34750,II34739,II34756,
    II34757,II34758,II34755,II34763,II34764,II34765,II34772,II34773,II34774,
    II34771,II34779,II34780,II34781,II34770,II34787,II34788,II34789,II34786,
    II34794,II34795,II34796,II34803,II34804,II34805,II34802,II34810,II34811,
    II34812,II34801,II34818,II34819,II34820,II34817,II34825,II34826,II34827,
    II34834,II34835,II34836,II34833,II34841,II34842,II34843,II34832,II34849,
    II34850,II34851,II34848,II34856,II34857,II34858,II34865,II34866,II34867,
    II34864,II34872,II34873,II34874,II34863,II34880,II34881,II34882,II34879,
    II34887,II34888,II34889,II34896,II34897,II34898,II34895,II34903,II34904,
    II34905,II34894,II34911,II34912,II34913,II34910,II34918,II34919,II34920,
    II34927,II34928,II34929,II34926,II34934,II34935,II34936,II34925,II34942,
    II34943,II34944,II34941,II34949,II34950,II34951,II34958,II34959,II34960,
    II34957,II34965,II34966,II34967,II34956,II34973,II34974,II34975,II34972,
    II34980,II34981,II34982,II34989,II34990,II34991,II34988,II34996,II34997,
    II34998,II34987,II35004,II35005,II35006,II35003,II35011,II35012,II35013,
    II35092,II35093,II35094,II35105,II35106,II35107,II35118,II35119,II35120,
    II35131,II35132,II35133,II35144,II35145,II35146,II35157,II35158,II35159,
    II35170,II35171,II35172,II35183,II35184,II35185,II35196,II35197,II35198,
    II35209,II35210,II35211,II35222,II35223,II35224,II35235,II35236,II35237,
    II35248,II35249,II35250,II35261,II35262,II35263,II35274,II35275,II35276,
    II35287,II35288,II35289,II35300,II35301,II35302,II35313,II35314,II35315,
    II35326,II35327,II35328,II35339,II35340,II35341,II35352,II35353,II35354,
    II35365,II35366,II35367,II35378,II35379,II35380,II35391,II35392,II35393,
    II35404,II35405,II35406,II35417,II35418,II35419,II35430,II35431,II35432,
    II35443,II35444,II35445,II35456,II35457,II35458,II35469,II35470,II35471,
    II35482,II35483,II35484,II35495,II35496,II35497,II35510,II35511,II35512,
    II35509,II35517,II35518,II35519,II35525,II35526,II35527,II35524,II35532,
    II35533,II35534,II35540,II35541,II35542,II35539,II35547,II35548,II35549,
    II35554,II35555,II35556,II35561,II35562,II35563,II35568,II35569,II35570,
    II35575,II35576,II35577,II35582,II35583,II35584,II35589,II35590,II35591,
    II35596,II35597,II35598,II35603,II35604,II35605,II35610,II35611,II35612,
    II35617,II35618,II35619,II35624,II35625,II35626,II35631,II35632,II35633,
    II35638,II35639,II35640,II35645,II35646,II35647,II35652,II35653,II35654,
    II35659,II35660,II35661,II35666,II35667,II35668,II35673,II35674,II35675,
    II35680,II35681,II35682,II35687,II35688,II35689,II35694,II35695,II35696,
    II35701,II35702,II35703,II35708,II35709,II35710,II35715,II35716,II35717,
    II35722,II35723,II35724,II35729,II35730,II35731,II35736,II35737,II35738,
    II35743,II35744,II35745,II35750,II35751,II35752;

  dff DFF_0(CK,WX485,WX484);
  dff DFF_1(CK,WX487,WX486);
  dff DFF_2(CK,WX489,WX488);
  dff DFF_3(CK,WX491,WX490);
  dff DFF_4(CK,WX493,WX492);
  dff DFF_5(CK,WX495,WX494);
  dff DFF_6(CK,WX497,WX496);
  dff DFF_7(CK,WX499,WX498);
  dff DFF_8(CK,WX501,WX500);
  dff DFF_9(CK,WX503,WX502);
  dff DFF_10(CK,WX505,WX504);
  dff DFF_11(CK,WX507,WX506);
  dff DFF_12(CK,WX509,WX508);
  dff DFF_13(CK,WX511,WX510);
  dff DFF_14(CK,WX513,WX512);
  dff DFF_15(CK,WX515,WX514);
  dff DFF_16(CK,WX517,WX516);
  dff DFF_17(CK,WX519,WX518);
  dff DFF_18(CK,WX521,WX520);
  dff DFF_19(CK,WX523,WX522);
  dff DFF_20(CK,WX525,WX524);
  dff DFF_21(CK,WX527,WX526);
  dff DFF_22(CK,WX529,WX528);
  dff DFF_23(CK,WX531,WX530);
  dff DFF_24(CK,WX533,WX532);
  dff DFF_25(CK,WX535,WX534);
  dff DFF_26(CK,WX537,WX536);
  dff DFF_27(CK,WX539,WX538);
  dff DFF_28(CK,WX541,WX540);
  dff DFF_29(CK,WX543,WX542);
  dff DFF_30(CK,WX545,WX544);
  dff DFF_31(CK,WX547,WX546);
  dff DFF_32(CK,WX645,WX644);
  dff DFF_33(CK,WX647,WX646);
  dff DFF_34(CK,WX649,WX648);
  dff DFF_35(CK,WX651,WX650);
  dff DFF_36(CK,WX653,WX652);
  dff DFF_37(CK,WX655,WX654);
  dff DFF_38(CK,WX657,WX656);
  dff DFF_39(CK,WX659,WX658);
  dff DFF_40(CK,WX661,WX660);
  dff DFF_41(CK,WX663,WX662);
  dff DFF_42(CK,WX665,WX664);
  dff DFF_43(CK,WX667,WX666);
  dff DFF_44(CK,WX669,WX668);
  dff DFF_45(CK,WX671,WX670);
  dff DFF_46(CK,WX673,WX672);
  dff DFF_47(CK,WX675,WX674);
  dff DFF_48(CK,WX677,WX676);
  dff DFF_49(CK,WX679,WX678);
  dff DFF_50(CK,WX681,WX680);
  dff DFF_51(CK,WX683,WX682);
  dff DFF_52(CK,WX685,WX684);
  dff DFF_53(CK,WX687,WX686);
  dff DFF_54(CK,WX689,WX688);
  dff DFF_55(CK,WX691,WX690);
  dff DFF_56(CK,WX693,WX692);
  dff DFF_57(CK,WX695,WX694);
  dff DFF_58(CK,WX697,WX696);
  dff DFF_59(CK,WX699,WX698);
  dff DFF_60(CK,WX701,WX700);
  dff DFF_61(CK,WX703,WX702);
  dff DFF_62(CK,WX705,WX704);
  dff DFF_63(CK,WX707,WX706);
  dff DFF_64(CK,WX709,WX708);
  dff DFF_65(CK,WX711,WX710);
  dff DFF_66(CK,WX713,WX712);
  dff DFF_67(CK,WX715,WX714);
  dff DFF_68(CK,WX717,WX716);
  dff DFF_69(CK,WX719,WX718);
  dff DFF_70(CK,WX721,WX720);
  dff DFF_71(CK,WX723,WX722);
  dff DFF_72(CK,WX725,WX724);
  dff DFF_73(CK,WX727,WX726);
  dff DFF_74(CK,WX729,WX728);
  dff DFF_75(CK,WX731,WX730);
  dff DFF_76(CK,WX733,WX732);
  dff DFF_77(CK,WX735,WX734);
  dff DFF_78(CK,WX737,WX736);
  dff DFF_79(CK,WX739,WX738);
  dff DFF_80(CK,WX741,WX740);
  dff DFF_81(CK,WX743,WX742);
  dff DFF_82(CK,WX745,WX744);
  dff DFF_83(CK,WX747,WX746);
  dff DFF_84(CK,WX749,WX748);
  dff DFF_85(CK,WX751,WX750);
  dff DFF_86(CK,WX753,WX752);
  dff DFF_87(CK,WX755,WX754);
  dff DFF_88(CK,WX757,WX756);
  dff DFF_89(CK,WX759,WX758);
  dff DFF_90(CK,WX761,WX760);
  dff DFF_91(CK,WX763,WX762);
  dff DFF_92(CK,WX765,WX764);
  dff DFF_93(CK,WX767,WX766);
  dff DFF_94(CK,WX769,WX768);
  dff DFF_95(CK,WX771,WX770);
  dff DFF_96(CK,WX773,WX772);
  dff DFF_97(CK,WX775,WX774);
  dff DFF_98(CK,WX777,WX776);
  dff DFF_99(CK,WX779,WX778);
  dff DFF_100(CK,WX781,WX780);
  dff DFF_101(CK,WX783,WX782);
  dff DFF_102(CK,WX785,WX784);
  dff DFF_103(CK,WX787,WX786);
  dff DFF_104(CK,WX789,WX788);
  dff DFF_105(CK,WX791,WX790);
  dff DFF_106(CK,WX793,WX792);
  dff DFF_107(CK,WX795,WX794);
  dff DFF_108(CK,WX797,WX796);
  dff DFF_109(CK,WX799,WX798);
  dff DFF_110(CK,WX801,WX800);
  dff DFF_111(CK,WX803,WX802);
  dff DFF_112(CK,WX805,WX804);
  dff DFF_113(CK,WX807,WX806);
  dff DFF_114(CK,WX809,WX808);
  dff DFF_115(CK,WX811,WX810);
  dff DFF_116(CK,WX813,WX812);
  dff DFF_117(CK,WX815,WX814);
  dff DFF_118(CK,WX817,WX816);
  dff DFF_119(CK,WX819,WX818);
  dff DFF_120(CK,WX821,WX820);
  dff DFF_121(CK,WX823,WX822);
  dff DFF_122(CK,WX825,WX824);
  dff DFF_123(CK,WX827,WX826);
  dff DFF_124(CK,WX829,WX828);
  dff DFF_125(CK,WX831,WX830);
  dff DFF_126(CK,WX833,WX832);
  dff DFF_127(CK,WX835,WX834);
  dff DFF_128(CK,WX837,WX836);
  dff DFF_129(CK,WX839,WX838);
  dff DFF_130(CK,WX841,WX840);
  dff DFF_131(CK,WX843,WX842);
  dff DFF_132(CK,WX845,WX844);
  dff DFF_133(CK,WX847,WX846);
  dff DFF_134(CK,WX849,WX848);
  dff DFF_135(CK,WX851,WX850);
  dff DFF_136(CK,WX853,WX852);
  dff DFF_137(CK,WX855,WX854);
  dff DFF_138(CK,WX857,WX856);
  dff DFF_139(CK,WX859,WX858);
  dff DFF_140(CK,WX861,WX860);
  dff DFF_141(CK,WX863,WX862);
  dff DFF_142(CK,WX865,WX864);
  dff DFF_143(CK,WX867,WX866);
  dff DFF_144(CK,WX869,WX868);
  dff DFF_145(CK,WX871,WX870);
  dff DFF_146(CK,WX873,WX872);
  dff DFF_147(CK,WX875,WX874);
  dff DFF_148(CK,WX877,WX876);
  dff DFF_149(CK,WX879,WX878);
  dff DFF_150(CK,WX881,WX880);
  dff DFF_151(CK,WX883,WX882);
  dff DFF_152(CK,WX885,WX884);
  dff DFF_153(CK,WX887,WX886);
  dff DFF_154(CK,WX889,WX888);
  dff DFF_155(CK,WX891,WX890);
  dff DFF_156(CK,WX893,WX892);
  dff DFF_157(CK,WX895,WX894);
  dff DFF_158(CK,WX897,WX896);
  dff DFF_159(CK,WX899,WX898);
  dff DFF_160(CK,CRC_OUT_9_0,WX1264);
  dff DFF_161(CK,CRC_OUT_9_1,WX1266);
  dff DFF_162(CK,CRC_OUT_9_2,WX1268);
  dff DFF_163(CK,CRC_OUT_9_3,WX1270);
  dff DFF_164(CK,CRC_OUT_9_4,WX1272);
  dff DFF_165(CK,CRC_OUT_9_5,WX1274);
  dff DFF_166(CK,CRC_OUT_9_6,WX1276);
  dff DFF_167(CK,CRC_OUT_9_7,WX1278);
  dff DFF_168(CK,CRC_OUT_9_8,WX1280);
  dff DFF_169(CK,CRC_OUT_9_9,WX1282);
  dff DFF_170(CK,CRC_OUT_9_10,WX1284);
  dff DFF_171(CK,CRC_OUT_9_11,WX1286);
  dff DFF_172(CK,CRC_OUT_9_12,WX1288);
  dff DFF_173(CK,CRC_OUT_9_13,WX1290);
  dff DFF_174(CK,CRC_OUT_9_14,WX1292);
  dff DFF_175(CK,CRC_OUT_9_15,WX1294);
  dff DFF_176(CK,CRC_OUT_9_16,WX1296);
  dff DFF_177(CK,CRC_OUT_9_17,WX1298);
  dff DFF_178(CK,CRC_OUT_9_18,WX1300);
  dff DFF_179(CK,CRC_OUT_9_19,WX1302);
  dff DFF_180(CK,CRC_OUT_9_20,WX1304);
  dff DFF_181(CK,CRC_OUT_9_21,WX1306);
  dff DFF_182(CK,CRC_OUT_9_22,WX1308);
  dff DFF_183(CK,CRC_OUT_9_23,WX1310);
  dff DFF_184(CK,CRC_OUT_9_24,WX1312);
  dff DFF_185(CK,CRC_OUT_9_25,WX1314);
  dff DFF_186(CK,CRC_OUT_9_26,WX1316);
  dff DFF_187(CK,CRC_OUT_9_27,WX1318);
  dff DFF_188(CK,CRC_OUT_9_28,WX1320);
  dff DFF_189(CK,CRC_OUT_9_29,WX1322);
  dff DFF_190(CK,CRC_OUT_9_30,WX1324);
  dff DFF_191(CK,CRC_OUT_9_31,WX1326);
  dff DFF_192(CK,WX1778,WX1777);
  dff DFF_193(CK,WX1780,WX1779);
  dff DFF_194(CK,WX1782,WX1781);
  dff DFF_195(CK,WX1784,WX1783);
  dff DFF_196(CK,WX1786,WX1785);
  dff DFF_197(CK,WX1788,WX1787);
  dff DFF_198(CK,WX1790,WX1789);
  dff DFF_199(CK,WX1792,WX1791);
  dff DFF_200(CK,WX1794,WX1793);
  dff DFF_201(CK,WX1796,WX1795);
  dff DFF_202(CK,WX1798,WX1797);
  dff DFF_203(CK,WX1800,WX1799);
  dff DFF_204(CK,WX1802,WX1801);
  dff DFF_205(CK,WX1804,WX1803);
  dff DFF_206(CK,WX1806,WX1805);
  dff DFF_207(CK,WX1808,WX1807);
  dff DFF_208(CK,WX1810,WX1809);
  dff DFF_209(CK,WX1812,WX1811);
  dff DFF_210(CK,WX1814,WX1813);
  dff DFF_211(CK,WX1816,WX1815);
  dff DFF_212(CK,WX1818,WX1817);
  dff DFF_213(CK,WX1820,WX1819);
  dff DFF_214(CK,WX1822,WX1821);
  dff DFF_215(CK,WX1824,WX1823);
  dff DFF_216(CK,WX1826,WX1825);
  dff DFF_217(CK,WX1828,WX1827);
  dff DFF_218(CK,WX1830,WX1829);
  dff DFF_219(CK,WX1832,WX1831);
  dff DFF_220(CK,WX1834,WX1833);
  dff DFF_221(CK,WX1836,WX1835);
  dff DFF_222(CK,WX1838,WX1837);
  dff DFF_223(CK,WX1840,WX1839);
  dff DFF_224(CK,WX1938,WX1937);
  dff DFF_225(CK,WX1940,WX1939);
  dff DFF_226(CK,WX1942,WX1941);
  dff DFF_227(CK,WX1944,WX1943);
  dff DFF_228(CK,WX1946,WX1945);
  dff DFF_229(CK,WX1948,WX1947);
  dff DFF_230(CK,WX1950,WX1949);
  dff DFF_231(CK,WX1952,WX1951);
  dff DFF_232(CK,WX1954,WX1953);
  dff DFF_233(CK,WX1956,WX1955);
  dff DFF_234(CK,WX1958,WX1957);
  dff DFF_235(CK,WX1960,WX1959);
  dff DFF_236(CK,WX1962,WX1961);
  dff DFF_237(CK,WX1964,WX1963);
  dff DFF_238(CK,WX1966,WX1965);
  dff DFF_239(CK,WX1968,WX1967);
  dff DFF_240(CK,WX1970,WX1969);
  dff DFF_241(CK,WX1972,WX1971);
  dff DFF_242(CK,WX1974,WX1973);
  dff DFF_243(CK,WX1976,WX1975);
  dff DFF_244(CK,WX1978,WX1977);
  dff DFF_245(CK,WX1980,WX1979);
  dff DFF_246(CK,WX1982,WX1981);
  dff DFF_247(CK,WX1984,WX1983);
  dff DFF_248(CK,WX1986,WX1985);
  dff DFF_249(CK,WX1988,WX1987);
  dff DFF_250(CK,WX1990,WX1989);
  dff DFF_251(CK,WX1992,WX1991);
  dff DFF_252(CK,WX1994,WX1993);
  dff DFF_253(CK,WX1996,WX1995);
  dff DFF_254(CK,WX1998,WX1997);
  dff DFF_255(CK,WX2000,WX1999);
  dff DFF_256(CK,WX2002,WX2001);
  dff DFF_257(CK,WX2004,WX2003);
  dff DFF_258(CK,WX2006,WX2005);
  dff DFF_259(CK,WX2008,WX2007);
  dff DFF_260(CK,WX2010,WX2009);
  dff DFF_261(CK,WX2012,WX2011);
  dff DFF_262(CK,WX2014,WX2013);
  dff DFF_263(CK,WX2016,WX2015);
  dff DFF_264(CK,WX2018,WX2017);
  dff DFF_265(CK,WX2020,WX2019);
  dff DFF_266(CK,WX2022,WX2021);
  dff DFF_267(CK,WX2024,WX2023);
  dff DFF_268(CK,WX2026,WX2025);
  dff DFF_269(CK,WX2028,WX2027);
  dff DFF_270(CK,WX2030,WX2029);
  dff DFF_271(CK,WX2032,WX2031);
  dff DFF_272(CK,WX2034,WX2033);
  dff DFF_273(CK,WX2036,WX2035);
  dff DFF_274(CK,WX2038,WX2037);
  dff DFF_275(CK,WX2040,WX2039);
  dff DFF_276(CK,WX2042,WX2041);
  dff DFF_277(CK,WX2044,WX2043);
  dff DFF_278(CK,WX2046,WX2045);
  dff DFF_279(CK,WX2048,WX2047);
  dff DFF_280(CK,WX2050,WX2049);
  dff DFF_281(CK,WX2052,WX2051);
  dff DFF_282(CK,WX2054,WX2053);
  dff DFF_283(CK,WX2056,WX2055);
  dff DFF_284(CK,WX2058,WX2057);
  dff DFF_285(CK,WX2060,WX2059);
  dff DFF_286(CK,WX2062,WX2061);
  dff DFF_287(CK,WX2064,WX2063);
  dff DFF_288(CK,WX2066,WX2065);
  dff DFF_289(CK,WX2068,WX2067);
  dff DFF_290(CK,WX2070,WX2069);
  dff DFF_291(CK,WX2072,WX2071);
  dff DFF_292(CK,WX2074,WX2073);
  dff DFF_293(CK,WX2076,WX2075);
  dff DFF_294(CK,WX2078,WX2077);
  dff DFF_295(CK,WX2080,WX2079);
  dff DFF_296(CK,WX2082,WX2081);
  dff DFF_297(CK,WX2084,WX2083);
  dff DFF_298(CK,WX2086,WX2085);
  dff DFF_299(CK,WX2088,WX2087);
  dff DFF_300(CK,WX2090,WX2089);
  dff DFF_301(CK,WX2092,WX2091);
  dff DFF_302(CK,WX2094,WX2093);
  dff DFF_303(CK,WX2096,WX2095);
  dff DFF_304(CK,WX2098,WX2097);
  dff DFF_305(CK,WX2100,WX2099);
  dff DFF_306(CK,WX2102,WX2101);
  dff DFF_307(CK,WX2104,WX2103);
  dff DFF_308(CK,WX2106,WX2105);
  dff DFF_309(CK,WX2108,WX2107);
  dff DFF_310(CK,WX2110,WX2109);
  dff DFF_311(CK,WX2112,WX2111);
  dff DFF_312(CK,WX2114,WX2113);
  dff DFF_313(CK,WX2116,WX2115);
  dff DFF_314(CK,WX2118,WX2117);
  dff DFF_315(CK,WX2120,WX2119);
  dff DFF_316(CK,WX2122,WX2121);
  dff DFF_317(CK,WX2124,WX2123);
  dff DFF_318(CK,WX2126,WX2125);
  dff DFF_319(CK,WX2128,WX2127);
  dff DFF_320(CK,WX2130,WX2129);
  dff DFF_321(CK,WX2132,WX2131);
  dff DFF_322(CK,WX2134,WX2133);
  dff DFF_323(CK,WX2136,WX2135);
  dff DFF_324(CK,WX2138,WX2137);
  dff DFF_325(CK,WX2140,WX2139);
  dff DFF_326(CK,WX2142,WX2141);
  dff DFF_327(CK,WX2144,WX2143);
  dff DFF_328(CK,WX2146,WX2145);
  dff DFF_329(CK,WX2148,WX2147);
  dff DFF_330(CK,WX2150,WX2149);
  dff DFF_331(CK,WX2152,WX2151);
  dff DFF_332(CK,WX2154,WX2153);
  dff DFF_333(CK,WX2156,WX2155);
  dff DFF_334(CK,WX2158,WX2157);
  dff DFF_335(CK,WX2160,WX2159);
  dff DFF_336(CK,WX2162,WX2161);
  dff DFF_337(CK,WX2164,WX2163);
  dff DFF_338(CK,WX2166,WX2165);
  dff DFF_339(CK,WX2168,WX2167);
  dff DFF_340(CK,WX2170,WX2169);
  dff DFF_341(CK,WX2172,WX2171);
  dff DFF_342(CK,WX2174,WX2173);
  dff DFF_343(CK,WX2176,WX2175);
  dff DFF_344(CK,WX2178,WX2177);
  dff DFF_345(CK,WX2180,WX2179);
  dff DFF_346(CK,WX2182,WX2181);
  dff DFF_347(CK,WX2184,WX2183);
  dff DFF_348(CK,WX2186,WX2185);
  dff DFF_349(CK,WX2188,WX2187);
  dff DFF_350(CK,WX2190,WX2189);
  dff DFF_351(CK,WX2192,WX2191);
  dff DFF_352(CK,CRC_OUT_8_0,WX2557);
  dff DFF_353(CK,CRC_OUT_8_1,WX2559);
  dff DFF_354(CK,CRC_OUT_8_2,WX2561);
  dff DFF_355(CK,CRC_OUT_8_3,WX2563);
  dff DFF_356(CK,CRC_OUT_8_4,WX2565);
  dff DFF_357(CK,CRC_OUT_8_5,WX2567);
  dff DFF_358(CK,CRC_OUT_8_6,WX2569);
  dff DFF_359(CK,CRC_OUT_8_7,WX2571);
  dff DFF_360(CK,CRC_OUT_8_8,WX2573);
  dff DFF_361(CK,CRC_OUT_8_9,WX2575);
  dff DFF_362(CK,CRC_OUT_8_10,WX2577);
  dff DFF_363(CK,CRC_OUT_8_11,WX2579);
  dff DFF_364(CK,CRC_OUT_8_12,WX2581);
  dff DFF_365(CK,CRC_OUT_8_13,WX2583);
  dff DFF_366(CK,CRC_OUT_8_14,WX2585);
  dff DFF_367(CK,CRC_OUT_8_15,WX2587);
  dff DFF_368(CK,CRC_OUT_8_16,WX2589);
  dff DFF_369(CK,CRC_OUT_8_17,WX2591);
  dff DFF_370(CK,CRC_OUT_8_18,WX2593);
  dff DFF_371(CK,CRC_OUT_8_19,WX2595);
  dff DFF_372(CK,CRC_OUT_8_20,WX2597);
  dff DFF_373(CK,CRC_OUT_8_21,WX2599);
  dff DFF_374(CK,CRC_OUT_8_22,WX2601);
  dff DFF_375(CK,CRC_OUT_8_23,WX2603);
  dff DFF_376(CK,CRC_OUT_8_24,WX2605);
  dff DFF_377(CK,CRC_OUT_8_25,WX2607);
  dff DFF_378(CK,CRC_OUT_8_26,WX2609);
  dff DFF_379(CK,CRC_OUT_8_27,WX2611);
  dff DFF_380(CK,CRC_OUT_8_28,WX2613);
  dff DFF_381(CK,CRC_OUT_8_29,WX2615);
  dff DFF_382(CK,CRC_OUT_8_30,WX2617);
  dff DFF_383(CK,CRC_OUT_8_31,WX2619);
  dff DFF_384(CK,WX3071,WX3070);
  dff DFF_385(CK,WX3073,WX3072);
  dff DFF_386(CK,WX3075,WX3074);
  dff DFF_387(CK,WX3077,WX3076);
  dff DFF_388(CK,WX3079,WX3078);
  dff DFF_389(CK,WX3081,WX3080);
  dff DFF_390(CK,WX3083,WX3082);
  dff DFF_391(CK,WX3085,WX3084);
  dff DFF_392(CK,WX3087,WX3086);
  dff DFF_393(CK,WX3089,WX3088);
  dff DFF_394(CK,WX3091,WX3090);
  dff DFF_395(CK,WX3093,WX3092);
  dff DFF_396(CK,WX3095,WX3094);
  dff DFF_397(CK,WX3097,WX3096);
  dff DFF_398(CK,WX3099,WX3098);
  dff DFF_399(CK,WX3101,WX3100);
  dff DFF_400(CK,WX3103,WX3102);
  dff DFF_401(CK,WX3105,WX3104);
  dff DFF_402(CK,WX3107,WX3106);
  dff DFF_403(CK,WX3109,WX3108);
  dff DFF_404(CK,WX3111,WX3110);
  dff DFF_405(CK,WX3113,WX3112);
  dff DFF_406(CK,WX3115,WX3114);
  dff DFF_407(CK,WX3117,WX3116);
  dff DFF_408(CK,WX3119,WX3118);
  dff DFF_409(CK,WX3121,WX3120);
  dff DFF_410(CK,WX3123,WX3122);
  dff DFF_411(CK,WX3125,WX3124);
  dff DFF_412(CK,WX3127,WX3126);
  dff DFF_413(CK,WX3129,WX3128);
  dff DFF_414(CK,WX3131,WX3130);
  dff DFF_415(CK,WX3133,WX3132);
  dff DFF_416(CK,WX3231,WX3230);
  dff DFF_417(CK,WX3233,WX3232);
  dff DFF_418(CK,WX3235,WX3234);
  dff DFF_419(CK,WX3237,WX3236);
  dff DFF_420(CK,WX3239,WX3238);
  dff DFF_421(CK,WX3241,WX3240);
  dff DFF_422(CK,WX3243,WX3242);
  dff DFF_423(CK,WX3245,WX3244);
  dff DFF_424(CK,WX3247,WX3246);
  dff DFF_425(CK,WX3249,WX3248);
  dff DFF_426(CK,WX3251,WX3250);
  dff DFF_427(CK,WX3253,WX3252);
  dff DFF_428(CK,WX3255,WX3254);
  dff DFF_429(CK,WX3257,WX3256);
  dff DFF_430(CK,WX3259,WX3258);
  dff DFF_431(CK,WX3261,WX3260);
  dff DFF_432(CK,WX3263,WX3262);
  dff DFF_433(CK,WX3265,WX3264);
  dff DFF_434(CK,WX3267,WX3266);
  dff DFF_435(CK,WX3269,WX3268);
  dff DFF_436(CK,WX3271,WX3270);
  dff DFF_437(CK,WX3273,WX3272);
  dff DFF_438(CK,WX3275,WX3274);
  dff DFF_439(CK,WX3277,WX3276);
  dff DFF_440(CK,WX3279,WX3278);
  dff DFF_441(CK,WX3281,WX3280);
  dff DFF_442(CK,WX3283,WX3282);
  dff DFF_443(CK,WX3285,WX3284);
  dff DFF_444(CK,WX3287,WX3286);
  dff DFF_445(CK,WX3289,WX3288);
  dff DFF_446(CK,WX3291,WX3290);
  dff DFF_447(CK,WX3293,WX3292);
  dff DFF_448(CK,WX3295,WX3294);
  dff DFF_449(CK,WX3297,WX3296);
  dff DFF_450(CK,WX3299,WX3298);
  dff DFF_451(CK,WX3301,WX3300);
  dff DFF_452(CK,WX3303,WX3302);
  dff DFF_453(CK,WX3305,WX3304);
  dff DFF_454(CK,WX3307,WX3306);
  dff DFF_455(CK,WX3309,WX3308);
  dff DFF_456(CK,WX3311,WX3310);
  dff DFF_457(CK,WX3313,WX3312);
  dff DFF_458(CK,WX3315,WX3314);
  dff DFF_459(CK,WX3317,WX3316);
  dff DFF_460(CK,WX3319,WX3318);
  dff DFF_461(CK,WX3321,WX3320);
  dff DFF_462(CK,WX3323,WX3322);
  dff DFF_463(CK,WX3325,WX3324);
  dff DFF_464(CK,WX3327,WX3326);
  dff DFF_465(CK,WX3329,WX3328);
  dff DFF_466(CK,WX3331,WX3330);
  dff DFF_467(CK,WX3333,WX3332);
  dff DFF_468(CK,WX3335,WX3334);
  dff DFF_469(CK,WX3337,WX3336);
  dff DFF_470(CK,WX3339,WX3338);
  dff DFF_471(CK,WX3341,WX3340);
  dff DFF_472(CK,WX3343,WX3342);
  dff DFF_473(CK,WX3345,WX3344);
  dff DFF_474(CK,WX3347,WX3346);
  dff DFF_475(CK,WX3349,WX3348);
  dff DFF_476(CK,WX3351,WX3350);
  dff DFF_477(CK,WX3353,WX3352);
  dff DFF_478(CK,WX3355,WX3354);
  dff DFF_479(CK,WX3357,WX3356);
  dff DFF_480(CK,WX3359,WX3358);
  dff DFF_481(CK,WX3361,WX3360);
  dff DFF_482(CK,WX3363,WX3362);
  dff DFF_483(CK,WX3365,WX3364);
  dff DFF_484(CK,WX3367,WX3366);
  dff DFF_485(CK,WX3369,WX3368);
  dff DFF_486(CK,WX3371,WX3370);
  dff DFF_487(CK,WX3373,WX3372);
  dff DFF_488(CK,WX3375,WX3374);
  dff DFF_489(CK,WX3377,WX3376);
  dff DFF_490(CK,WX3379,WX3378);
  dff DFF_491(CK,WX3381,WX3380);
  dff DFF_492(CK,WX3383,WX3382);
  dff DFF_493(CK,WX3385,WX3384);
  dff DFF_494(CK,WX3387,WX3386);
  dff DFF_495(CK,WX3389,WX3388);
  dff DFF_496(CK,WX3391,WX3390);
  dff DFF_497(CK,WX3393,WX3392);
  dff DFF_498(CK,WX3395,WX3394);
  dff DFF_499(CK,WX3397,WX3396);
  dff DFF_500(CK,WX3399,WX3398);
  dff DFF_501(CK,WX3401,WX3400);
  dff DFF_502(CK,WX3403,WX3402);
  dff DFF_503(CK,WX3405,WX3404);
  dff DFF_504(CK,WX3407,WX3406);
  dff DFF_505(CK,WX3409,WX3408);
  dff DFF_506(CK,WX3411,WX3410);
  dff DFF_507(CK,WX3413,WX3412);
  dff DFF_508(CK,WX3415,WX3414);
  dff DFF_509(CK,WX3417,WX3416);
  dff DFF_510(CK,WX3419,WX3418);
  dff DFF_511(CK,WX3421,WX3420);
  dff DFF_512(CK,WX3423,WX3422);
  dff DFF_513(CK,WX3425,WX3424);
  dff DFF_514(CK,WX3427,WX3426);
  dff DFF_515(CK,WX3429,WX3428);
  dff DFF_516(CK,WX3431,WX3430);
  dff DFF_517(CK,WX3433,WX3432);
  dff DFF_518(CK,WX3435,WX3434);
  dff DFF_519(CK,WX3437,WX3436);
  dff DFF_520(CK,WX3439,WX3438);
  dff DFF_521(CK,WX3441,WX3440);
  dff DFF_522(CK,WX3443,WX3442);
  dff DFF_523(CK,WX3445,WX3444);
  dff DFF_524(CK,WX3447,WX3446);
  dff DFF_525(CK,WX3449,WX3448);
  dff DFF_526(CK,WX3451,WX3450);
  dff DFF_527(CK,WX3453,WX3452);
  dff DFF_528(CK,WX3455,WX3454);
  dff DFF_529(CK,WX3457,WX3456);
  dff DFF_530(CK,WX3459,WX3458);
  dff DFF_531(CK,WX3461,WX3460);
  dff DFF_532(CK,WX3463,WX3462);
  dff DFF_533(CK,WX3465,WX3464);
  dff DFF_534(CK,WX3467,WX3466);
  dff DFF_535(CK,WX3469,WX3468);
  dff DFF_536(CK,WX3471,WX3470);
  dff DFF_537(CK,WX3473,WX3472);
  dff DFF_538(CK,WX3475,WX3474);
  dff DFF_539(CK,WX3477,WX3476);
  dff DFF_540(CK,WX3479,WX3478);
  dff DFF_541(CK,WX3481,WX3480);
  dff DFF_542(CK,WX3483,WX3482);
  dff DFF_543(CK,WX3485,WX3484);
  dff DFF_544(CK,CRC_OUT_7_0,WX3850);
  dff DFF_545(CK,CRC_OUT_7_1,WX3852);
  dff DFF_546(CK,CRC_OUT_7_2,WX3854);
  dff DFF_547(CK,CRC_OUT_7_3,WX3856);
  dff DFF_548(CK,CRC_OUT_7_4,WX3858);
  dff DFF_549(CK,CRC_OUT_7_5,WX3860);
  dff DFF_550(CK,CRC_OUT_7_6,WX3862);
  dff DFF_551(CK,CRC_OUT_7_7,WX3864);
  dff DFF_552(CK,CRC_OUT_7_8,WX3866);
  dff DFF_553(CK,CRC_OUT_7_9,WX3868);
  dff DFF_554(CK,CRC_OUT_7_10,WX3870);
  dff DFF_555(CK,CRC_OUT_7_11,WX3872);
  dff DFF_556(CK,CRC_OUT_7_12,WX3874);
  dff DFF_557(CK,CRC_OUT_7_13,WX3876);
  dff DFF_558(CK,CRC_OUT_7_14,WX3878);
  dff DFF_559(CK,CRC_OUT_7_15,WX3880);
  dff DFF_560(CK,CRC_OUT_7_16,WX3882);
  dff DFF_561(CK,CRC_OUT_7_17,WX3884);
  dff DFF_562(CK,CRC_OUT_7_18,WX3886);
  dff DFF_563(CK,CRC_OUT_7_19,WX3888);
  dff DFF_564(CK,CRC_OUT_7_20,WX3890);
  dff DFF_565(CK,CRC_OUT_7_21,WX3892);
  dff DFF_566(CK,CRC_OUT_7_22,WX3894);
  dff DFF_567(CK,CRC_OUT_7_23,WX3896);
  dff DFF_568(CK,CRC_OUT_7_24,WX3898);
  dff DFF_569(CK,CRC_OUT_7_25,WX3900);
  dff DFF_570(CK,CRC_OUT_7_26,WX3902);
  dff DFF_571(CK,CRC_OUT_7_27,WX3904);
  dff DFF_572(CK,CRC_OUT_7_28,WX3906);
  dff DFF_573(CK,CRC_OUT_7_29,WX3908);
  dff DFF_574(CK,CRC_OUT_7_30,WX3910);
  dff DFF_575(CK,CRC_OUT_7_31,WX3912);
  dff DFF_576(CK,WX4364,WX4363);
  dff DFF_577(CK,WX4366,WX4365);
  dff DFF_578(CK,WX4368,WX4367);
  dff DFF_579(CK,WX4370,WX4369);
  dff DFF_580(CK,WX4372,WX4371);
  dff DFF_581(CK,WX4374,WX4373);
  dff DFF_582(CK,WX4376,WX4375);
  dff DFF_583(CK,WX4378,WX4377);
  dff DFF_584(CK,WX4380,WX4379);
  dff DFF_585(CK,WX4382,WX4381);
  dff DFF_586(CK,WX4384,WX4383);
  dff DFF_587(CK,WX4386,WX4385);
  dff DFF_588(CK,WX4388,WX4387);
  dff DFF_589(CK,WX4390,WX4389);
  dff DFF_590(CK,WX4392,WX4391);
  dff DFF_591(CK,WX4394,WX4393);
  dff DFF_592(CK,WX4396,WX4395);
  dff DFF_593(CK,WX4398,WX4397);
  dff DFF_594(CK,WX4400,WX4399);
  dff DFF_595(CK,WX4402,WX4401);
  dff DFF_596(CK,WX4404,WX4403);
  dff DFF_597(CK,WX4406,WX4405);
  dff DFF_598(CK,WX4408,WX4407);
  dff DFF_599(CK,WX4410,WX4409);
  dff DFF_600(CK,WX4412,WX4411);
  dff DFF_601(CK,WX4414,WX4413);
  dff DFF_602(CK,WX4416,WX4415);
  dff DFF_603(CK,WX4418,WX4417);
  dff DFF_604(CK,WX4420,WX4419);
  dff DFF_605(CK,WX4422,WX4421);
  dff DFF_606(CK,WX4424,WX4423);
  dff DFF_607(CK,WX4426,WX4425);
  dff DFF_608(CK,WX4524,WX4523);
  dff DFF_609(CK,WX4526,WX4525);
  dff DFF_610(CK,WX4528,WX4527);
  dff DFF_611(CK,WX4530,WX4529);
  dff DFF_612(CK,WX4532,WX4531);
  dff DFF_613(CK,WX4534,WX4533);
  dff DFF_614(CK,WX4536,WX4535);
  dff DFF_615(CK,WX4538,WX4537);
  dff DFF_616(CK,WX4540,WX4539);
  dff DFF_617(CK,WX4542,WX4541);
  dff DFF_618(CK,WX4544,WX4543);
  dff DFF_619(CK,WX4546,WX4545);
  dff DFF_620(CK,WX4548,WX4547);
  dff DFF_621(CK,WX4550,WX4549);
  dff DFF_622(CK,WX4552,WX4551);
  dff DFF_623(CK,WX4554,WX4553);
  dff DFF_624(CK,WX4556,WX4555);
  dff DFF_625(CK,WX4558,WX4557);
  dff DFF_626(CK,WX4560,WX4559);
  dff DFF_627(CK,WX4562,WX4561);
  dff DFF_628(CK,WX4564,WX4563);
  dff DFF_629(CK,WX4566,WX4565);
  dff DFF_630(CK,WX4568,WX4567);
  dff DFF_631(CK,WX4570,WX4569);
  dff DFF_632(CK,WX4572,WX4571);
  dff DFF_633(CK,WX4574,WX4573);
  dff DFF_634(CK,WX4576,WX4575);
  dff DFF_635(CK,WX4578,WX4577);
  dff DFF_636(CK,WX4580,WX4579);
  dff DFF_637(CK,WX4582,WX4581);
  dff DFF_638(CK,WX4584,WX4583);
  dff DFF_639(CK,WX4586,WX4585);
  dff DFF_640(CK,WX4588,WX4587);
  dff DFF_641(CK,WX4590,WX4589);
  dff DFF_642(CK,WX4592,WX4591);
  dff DFF_643(CK,WX4594,WX4593);
  dff DFF_644(CK,WX4596,WX4595);
  dff DFF_645(CK,WX4598,WX4597);
  dff DFF_646(CK,WX4600,WX4599);
  dff DFF_647(CK,WX4602,WX4601);
  dff DFF_648(CK,WX4604,WX4603);
  dff DFF_649(CK,WX4606,WX4605);
  dff DFF_650(CK,WX4608,WX4607);
  dff DFF_651(CK,WX4610,WX4609);
  dff DFF_652(CK,WX4612,WX4611);
  dff DFF_653(CK,WX4614,WX4613);
  dff DFF_654(CK,WX4616,WX4615);
  dff DFF_655(CK,WX4618,WX4617);
  dff DFF_656(CK,WX4620,WX4619);
  dff DFF_657(CK,WX4622,WX4621);
  dff DFF_658(CK,WX4624,WX4623);
  dff DFF_659(CK,WX4626,WX4625);
  dff DFF_660(CK,WX4628,WX4627);
  dff DFF_661(CK,WX4630,WX4629);
  dff DFF_662(CK,WX4632,WX4631);
  dff DFF_663(CK,WX4634,WX4633);
  dff DFF_664(CK,WX4636,WX4635);
  dff DFF_665(CK,WX4638,WX4637);
  dff DFF_666(CK,WX4640,WX4639);
  dff DFF_667(CK,WX4642,WX4641);
  dff DFF_668(CK,WX4644,WX4643);
  dff DFF_669(CK,WX4646,WX4645);
  dff DFF_670(CK,WX4648,WX4647);
  dff DFF_671(CK,WX4650,WX4649);
  dff DFF_672(CK,WX4652,WX4651);
  dff DFF_673(CK,WX4654,WX4653);
  dff DFF_674(CK,WX4656,WX4655);
  dff DFF_675(CK,WX4658,WX4657);
  dff DFF_676(CK,WX4660,WX4659);
  dff DFF_677(CK,WX4662,WX4661);
  dff DFF_678(CK,WX4664,WX4663);
  dff DFF_679(CK,WX4666,WX4665);
  dff DFF_680(CK,WX4668,WX4667);
  dff DFF_681(CK,WX4670,WX4669);
  dff DFF_682(CK,WX4672,WX4671);
  dff DFF_683(CK,WX4674,WX4673);
  dff DFF_684(CK,WX4676,WX4675);
  dff DFF_685(CK,WX4678,WX4677);
  dff DFF_686(CK,WX4680,WX4679);
  dff DFF_687(CK,WX4682,WX4681);
  dff DFF_688(CK,WX4684,WX4683);
  dff DFF_689(CK,WX4686,WX4685);
  dff DFF_690(CK,WX4688,WX4687);
  dff DFF_691(CK,WX4690,WX4689);
  dff DFF_692(CK,WX4692,WX4691);
  dff DFF_693(CK,WX4694,WX4693);
  dff DFF_694(CK,WX4696,WX4695);
  dff DFF_695(CK,WX4698,WX4697);
  dff DFF_696(CK,WX4700,WX4699);
  dff DFF_697(CK,WX4702,WX4701);
  dff DFF_698(CK,WX4704,WX4703);
  dff DFF_699(CK,WX4706,WX4705);
  dff DFF_700(CK,WX4708,WX4707);
  dff DFF_701(CK,WX4710,WX4709);
  dff DFF_702(CK,WX4712,WX4711);
  dff DFF_703(CK,WX4714,WX4713);
  dff DFF_704(CK,WX4716,WX4715);
  dff DFF_705(CK,WX4718,WX4717);
  dff DFF_706(CK,WX4720,WX4719);
  dff DFF_707(CK,WX4722,WX4721);
  dff DFF_708(CK,WX4724,WX4723);
  dff DFF_709(CK,WX4726,WX4725);
  dff DFF_710(CK,WX4728,WX4727);
  dff DFF_711(CK,WX4730,WX4729);
  dff DFF_712(CK,WX4732,WX4731);
  dff DFF_713(CK,WX4734,WX4733);
  dff DFF_714(CK,WX4736,WX4735);
  dff DFF_715(CK,WX4738,WX4737);
  dff DFF_716(CK,WX4740,WX4739);
  dff DFF_717(CK,WX4742,WX4741);
  dff DFF_718(CK,WX4744,WX4743);
  dff DFF_719(CK,WX4746,WX4745);
  dff DFF_720(CK,WX4748,WX4747);
  dff DFF_721(CK,WX4750,WX4749);
  dff DFF_722(CK,WX4752,WX4751);
  dff DFF_723(CK,WX4754,WX4753);
  dff DFF_724(CK,WX4756,WX4755);
  dff DFF_725(CK,WX4758,WX4757);
  dff DFF_726(CK,WX4760,WX4759);
  dff DFF_727(CK,WX4762,WX4761);
  dff DFF_728(CK,WX4764,WX4763);
  dff DFF_729(CK,WX4766,WX4765);
  dff DFF_730(CK,WX4768,WX4767);
  dff DFF_731(CK,WX4770,WX4769);
  dff DFF_732(CK,WX4772,WX4771);
  dff DFF_733(CK,WX4774,WX4773);
  dff DFF_734(CK,WX4776,WX4775);
  dff DFF_735(CK,WX4778,WX4777);
  dff DFF_736(CK,CRC_OUT_6_0,WX5143);
  dff DFF_737(CK,CRC_OUT_6_1,WX5145);
  dff DFF_738(CK,CRC_OUT_6_2,WX5147);
  dff DFF_739(CK,CRC_OUT_6_3,WX5149);
  dff DFF_740(CK,CRC_OUT_6_4,WX5151);
  dff DFF_741(CK,CRC_OUT_6_5,WX5153);
  dff DFF_742(CK,CRC_OUT_6_6,WX5155);
  dff DFF_743(CK,CRC_OUT_6_7,WX5157);
  dff DFF_744(CK,CRC_OUT_6_8,WX5159);
  dff DFF_745(CK,CRC_OUT_6_9,WX5161);
  dff DFF_746(CK,CRC_OUT_6_10,WX5163);
  dff DFF_747(CK,CRC_OUT_6_11,WX5165);
  dff DFF_748(CK,CRC_OUT_6_12,WX5167);
  dff DFF_749(CK,CRC_OUT_6_13,WX5169);
  dff DFF_750(CK,CRC_OUT_6_14,WX5171);
  dff DFF_751(CK,CRC_OUT_6_15,WX5173);
  dff DFF_752(CK,CRC_OUT_6_16,WX5175);
  dff DFF_753(CK,CRC_OUT_6_17,WX5177);
  dff DFF_754(CK,CRC_OUT_6_18,WX5179);
  dff DFF_755(CK,CRC_OUT_6_19,WX5181);
  dff DFF_756(CK,CRC_OUT_6_20,WX5183);
  dff DFF_757(CK,CRC_OUT_6_21,WX5185);
  dff DFF_758(CK,CRC_OUT_6_22,WX5187);
  dff DFF_759(CK,CRC_OUT_6_23,WX5189);
  dff DFF_760(CK,CRC_OUT_6_24,WX5191);
  dff DFF_761(CK,CRC_OUT_6_25,WX5193);
  dff DFF_762(CK,CRC_OUT_6_26,WX5195);
  dff DFF_763(CK,CRC_OUT_6_27,WX5197);
  dff DFF_764(CK,CRC_OUT_6_28,WX5199);
  dff DFF_765(CK,CRC_OUT_6_29,WX5201);
  dff DFF_766(CK,CRC_OUT_6_30,WX5203);
  dff DFF_767(CK,CRC_OUT_6_31,WX5205);
  dff DFF_768(CK,WX5657,WX5656);
  dff DFF_769(CK,WX5659,WX5658);
  dff DFF_770(CK,WX5661,WX5660);
  dff DFF_771(CK,WX5663,WX5662);
  dff DFF_772(CK,WX5665,WX5664);
  dff DFF_773(CK,WX5667,WX5666);
  dff DFF_774(CK,WX5669,WX5668);
  dff DFF_775(CK,WX5671,WX5670);
  dff DFF_776(CK,WX5673,WX5672);
  dff DFF_777(CK,WX5675,WX5674);
  dff DFF_778(CK,WX5677,WX5676);
  dff DFF_779(CK,WX5679,WX5678);
  dff DFF_780(CK,WX5681,WX5680);
  dff DFF_781(CK,WX5683,WX5682);
  dff DFF_782(CK,WX5685,WX5684);
  dff DFF_783(CK,WX5687,WX5686);
  dff DFF_784(CK,WX5689,WX5688);
  dff DFF_785(CK,WX5691,WX5690);
  dff DFF_786(CK,WX5693,WX5692);
  dff DFF_787(CK,WX5695,WX5694);
  dff DFF_788(CK,WX5697,WX5696);
  dff DFF_789(CK,WX5699,WX5698);
  dff DFF_790(CK,WX5701,WX5700);
  dff DFF_791(CK,WX5703,WX5702);
  dff DFF_792(CK,WX5705,WX5704);
  dff DFF_793(CK,WX5707,WX5706);
  dff DFF_794(CK,WX5709,WX5708);
  dff DFF_795(CK,WX5711,WX5710);
  dff DFF_796(CK,WX5713,WX5712);
  dff DFF_797(CK,WX5715,WX5714);
  dff DFF_798(CK,WX5717,WX5716);
  dff DFF_799(CK,WX5719,WX5718);
  dff DFF_800(CK,WX5817,WX5816);
  dff DFF_801(CK,WX5819,WX5818);
  dff DFF_802(CK,WX5821,WX5820);
  dff DFF_803(CK,WX5823,WX5822);
  dff DFF_804(CK,WX5825,WX5824);
  dff DFF_805(CK,WX5827,WX5826);
  dff DFF_806(CK,WX5829,WX5828);
  dff DFF_807(CK,WX5831,WX5830);
  dff DFF_808(CK,WX5833,WX5832);
  dff DFF_809(CK,WX5835,WX5834);
  dff DFF_810(CK,WX5837,WX5836);
  dff DFF_811(CK,WX5839,WX5838);
  dff DFF_812(CK,WX5841,WX5840);
  dff DFF_813(CK,WX5843,WX5842);
  dff DFF_814(CK,WX5845,WX5844);
  dff DFF_815(CK,WX5847,WX5846);
  dff DFF_816(CK,WX5849,WX5848);
  dff DFF_817(CK,WX5851,WX5850);
  dff DFF_818(CK,WX5853,WX5852);
  dff DFF_819(CK,WX5855,WX5854);
  dff DFF_820(CK,WX5857,WX5856);
  dff DFF_821(CK,WX5859,WX5858);
  dff DFF_822(CK,WX5861,WX5860);
  dff DFF_823(CK,WX5863,WX5862);
  dff DFF_824(CK,WX5865,WX5864);
  dff DFF_825(CK,WX5867,WX5866);
  dff DFF_826(CK,WX5869,WX5868);
  dff DFF_827(CK,WX5871,WX5870);
  dff DFF_828(CK,WX5873,WX5872);
  dff DFF_829(CK,WX5875,WX5874);
  dff DFF_830(CK,WX5877,WX5876);
  dff DFF_831(CK,WX5879,WX5878);
  dff DFF_832(CK,WX5881,WX5880);
  dff DFF_833(CK,WX5883,WX5882);
  dff DFF_834(CK,WX5885,WX5884);
  dff DFF_835(CK,WX5887,WX5886);
  dff DFF_836(CK,WX5889,WX5888);
  dff DFF_837(CK,WX5891,WX5890);
  dff DFF_838(CK,WX5893,WX5892);
  dff DFF_839(CK,WX5895,WX5894);
  dff DFF_840(CK,WX5897,WX5896);
  dff DFF_841(CK,WX5899,WX5898);
  dff DFF_842(CK,WX5901,WX5900);
  dff DFF_843(CK,WX5903,WX5902);
  dff DFF_844(CK,WX5905,WX5904);
  dff DFF_845(CK,WX5907,WX5906);
  dff DFF_846(CK,WX5909,WX5908);
  dff DFF_847(CK,WX5911,WX5910);
  dff DFF_848(CK,WX5913,WX5912);
  dff DFF_849(CK,WX5915,WX5914);
  dff DFF_850(CK,WX5917,WX5916);
  dff DFF_851(CK,WX5919,WX5918);
  dff DFF_852(CK,WX5921,WX5920);
  dff DFF_853(CK,WX5923,WX5922);
  dff DFF_854(CK,WX5925,WX5924);
  dff DFF_855(CK,WX5927,WX5926);
  dff DFF_856(CK,WX5929,WX5928);
  dff DFF_857(CK,WX5931,WX5930);
  dff DFF_858(CK,WX5933,WX5932);
  dff DFF_859(CK,WX5935,WX5934);
  dff DFF_860(CK,WX5937,WX5936);
  dff DFF_861(CK,WX5939,WX5938);
  dff DFF_862(CK,WX5941,WX5940);
  dff DFF_863(CK,WX5943,WX5942);
  dff DFF_864(CK,WX5945,WX5944);
  dff DFF_865(CK,WX5947,WX5946);
  dff DFF_866(CK,WX5949,WX5948);
  dff DFF_867(CK,WX5951,WX5950);
  dff DFF_868(CK,WX5953,WX5952);
  dff DFF_869(CK,WX5955,WX5954);
  dff DFF_870(CK,WX5957,WX5956);
  dff DFF_871(CK,WX5959,WX5958);
  dff DFF_872(CK,WX5961,WX5960);
  dff DFF_873(CK,WX5963,WX5962);
  dff DFF_874(CK,WX5965,WX5964);
  dff DFF_875(CK,WX5967,WX5966);
  dff DFF_876(CK,WX5969,WX5968);
  dff DFF_877(CK,WX5971,WX5970);
  dff DFF_878(CK,WX5973,WX5972);
  dff DFF_879(CK,WX5975,WX5974);
  dff DFF_880(CK,WX5977,WX5976);
  dff DFF_881(CK,WX5979,WX5978);
  dff DFF_882(CK,WX5981,WX5980);
  dff DFF_883(CK,WX5983,WX5982);
  dff DFF_884(CK,WX5985,WX5984);
  dff DFF_885(CK,WX5987,WX5986);
  dff DFF_886(CK,WX5989,WX5988);
  dff DFF_887(CK,WX5991,WX5990);
  dff DFF_888(CK,WX5993,WX5992);
  dff DFF_889(CK,WX5995,WX5994);
  dff DFF_890(CK,WX5997,WX5996);
  dff DFF_891(CK,WX5999,WX5998);
  dff DFF_892(CK,WX6001,WX6000);
  dff DFF_893(CK,WX6003,WX6002);
  dff DFF_894(CK,WX6005,WX6004);
  dff DFF_895(CK,WX6007,WX6006);
  dff DFF_896(CK,WX6009,WX6008);
  dff DFF_897(CK,WX6011,WX6010);
  dff DFF_898(CK,WX6013,WX6012);
  dff DFF_899(CK,WX6015,WX6014);
  dff DFF_900(CK,WX6017,WX6016);
  dff DFF_901(CK,WX6019,WX6018);
  dff DFF_902(CK,WX6021,WX6020);
  dff DFF_903(CK,WX6023,WX6022);
  dff DFF_904(CK,WX6025,WX6024);
  dff DFF_905(CK,WX6027,WX6026);
  dff DFF_906(CK,WX6029,WX6028);
  dff DFF_907(CK,WX6031,WX6030);
  dff DFF_908(CK,WX6033,WX6032);
  dff DFF_909(CK,WX6035,WX6034);
  dff DFF_910(CK,WX6037,WX6036);
  dff DFF_911(CK,WX6039,WX6038);
  dff DFF_912(CK,WX6041,WX6040);
  dff DFF_913(CK,WX6043,WX6042);
  dff DFF_914(CK,WX6045,WX6044);
  dff DFF_915(CK,WX6047,WX6046);
  dff DFF_916(CK,WX6049,WX6048);
  dff DFF_917(CK,WX6051,WX6050);
  dff DFF_918(CK,WX6053,WX6052);
  dff DFF_919(CK,WX6055,WX6054);
  dff DFF_920(CK,WX6057,WX6056);
  dff DFF_921(CK,WX6059,WX6058);
  dff DFF_922(CK,WX6061,WX6060);
  dff DFF_923(CK,WX6063,WX6062);
  dff DFF_924(CK,WX6065,WX6064);
  dff DFF_925(CK,WX6067,WX6066);
  dff DFF_926(CK,WX6069,WX6068);
  dff DFF_927(CK,WX6071,WX6070);
  dff DFF_928(CK,CRC_OUT_5_0,WX6436);
  dff DFF_929(CK,CRC_OUT_5_1,WX6438);
  dff DFF_930(CK,CRC_OUT_5_2,WX6440);
  dff DFF_931(CK,CRC_OUT_5_3,WX6442);
  dff DFF_932(CK,CRC_OUT_5_4,WX6444);
  dff DFF_933(CK,CRC_OUT_5_5,WX6446);
  dff DFF_934(CK,CRC_OUT_5_6,WX6448);
  dff DFF_935(CK,CRC_OUT_5_7,WX6450);
  dff DFF_936(CK,CRC_OUT_5_8,WX6452);
  dff DFF_937(CK,CRC_OUT_5_9,WX6454);
  dff DFF_938(CK,CRC_OUT_5_10,WX6456);
  dff DFF_939(CK,CRC_OUT_5_11,WX6458);
  dff DFF_940(CK,CRC_OUT_5_12,WX6460);
  dff DFF_941(CK,CRC_OUT_5_13,WX6462);
  dff DFF_942(CK,CRC_OUT_5_14,WX6464);
  dff DFF_943(CK,CRC_OUT_5_15,WX6466);
  dff DFF_944(CK,CRC_OUT_5_16,WX6468);
  dff DFF_945(CK,CRC_OUT_5_17,WX6470);
  dff DFF_946(CK,CRC_OUT_5_18,WX6472);
  dff DFF_947(CK,CRC_OUT_5_19,WX6474);
  dff DFF_948(CK,CRC_OUT_5_20,WX6476);
  dff DFF_949(CK,CRC_OUT_5_21,WX6478);
  dff DFF_950(CK,CRC_OUT_5_22,WX6480);
  dff DFF_951(CK,CRC_OUT_5_23,WX6482);
  dff DFF_952(CK,CRC_OUT_5_24,WX6484);
  dff DFF_953(CK,CRC_OUT_5_25,WX6486);
  dff DFF_954(CK,CRC_OUT_5_26,WX6488);
  dff DFF_955(CK,CRC_OUT_5_27,WX6490);
  dff DFF_956(CK,CRC_OUT_5_28,WX6492);
  dff DFF_957(CK,CRC_OUT_5_29,WX6494);
  dff DFF_958(CK,CRC_OUT_5_30,WX6496);
  dff DFF_959(CK,CRC_OUT_5_31,WX6498);
  dff DFF_960(CK,WX6950,WX6949);
  dff DFF_961(CK,WX6952,WX6951);
  dff DFF_962(CK,WX6954,WX6953);
  dff DFF_963(CK,WX6956,WX6955);
  dff DFF_964(CK,WX6958,WX6957);
  dff DFF_965(CK,WX6960,WX6959);
  dff DFF_966(CK,WX6962,WX6961);
  dff DFF_967(CK,WX6964,WX6963);
  dff DFF_968(CK,WX6966,WX6965);
  dff DFF_969(CK,WX6968,WX6967);
  dff DFF_970(CK,WX6970,WX6969);
  dff DFF_971(CK,WX6972,WX6971);
  dff DFF_972(CK,WX6974,WX6973);
  dff DFF_973(CK,WX6976,WX6975);
  dff DFF_974(CK,WX6978,WX6977);
  dff DFF_975(CK,WX6980,WX6979);
  dff DFF_976(CK,WX6982,WX6981);
  dff DFF_977(CK,WX6984,WX6983);
  dff DFF_978(CK,WX6986,WX6985);
  dff DFF_979(CK,WX6988,WX6987);
  dff DFF_980(CK,WX6990,WX6989);
  dff DFF_981(CK,WX6992,WX6991);
  dff DFF_982(CK,WX6994,WX6993);
  dff DFF_983(CK,WX6996,WX6995);
  dff DFF_984(CK,WX6998,WX6997);
  dff DFF_985(CK,WX7000,WX6999);
  dff DFF_986(CK,WX7002,WX7001);
  dff DFF_987(CK,WX7004,WX7003);
  dff DFF_988(CK,WX7006,WX7005);
  dff DFF_989(CK,WX7008,WX7007);
  dff DFF_990(CK,WX7010,WX7009);
  dff DFF_991(CK,WX7012,WX7011);
  dff DFF_992(CK,WX7110,WX7109);
  dff DFF_993(CK,WX7112,WX7111);
  dff DFF_994(CK,WX7114,WX7113);
  dff DFF_995(CK,WX7116,WX7115);
  dff DFF_996(CK,WX7118,WX7117);
  dff DFF_997(CK,WX7120,WX7119);
  dff DFF_998(CK,WX7122,WX7121);
  dff DFF_999(CK,WX7124,WX7123);
  dff DFF_1000(CK,WX7126,WX7125);
  dff DFF_1001(CK,WX7128,WX7127);
  dff DFF_1002(CK,WX7130,WX7129);
  dff DFF_1003(CK,WX7132,WX7131);
  dff DFF_1004(CK,WX7134,WX7133);
  dff DFF_1005(CK,WX7136,WX7135);
  dff DFF_1006(CK,WX7138,WX7137);
  dff DFF_1007(CK,WX7140,WX7139);
  dff DFF_1008(CK,WX7142,WX7141);
  dff DFF_1009(CK,WX7144,WX7143);
  dff DFF_1010(CK,WX7146,WX7145);
  dff DFF_1011(CK,WX7148,WX7147);
  dff DFF_1012(CK,WX7150,WX7149);
  dff DFF_1013(CK,WX7152,WX7151);
  dff DFF_1014(CK,WX7154,WX7153);
  dff DFF_1015(CK,WX7156,WX7155);
  dff DFF_1016(CK,WX7158,WX7157);
  dff DFF_1017(CK,WX7160,WX7159);
  dff DFF_1018(CK,WX7162,WX7161);
  dff DFF_1019(CK,WX7164,WX7163);
  dff DFF_1020(CK,WX7166,WX7165);
  dff DFF_1021(CK,WX7168,WX7167);
  dff DFF_1022(CK,WX7170,WX7169);
  dff DFF_1023(CK,WX7172,WX7171);
  dff DFF_1024(CK,WX7174,WX7173);
  dff DFF_1025(CK,WX7176,WX7175);
  dff DFF_1026(CK,WX7178,WX7177);
  dff DFF_1027(CK,WX7180,WX7179);
  dff DFF_1028(CK,WX7182,WX7181);
  dff DFF_1029(CK,WX7184,WX7183);
  dff DFF_1030(CK,WX7186,WX7185);
  dff DFF_1031(CK,WX7188,WX7187);
  dff DFF_1032(CK,WX7190,WX7189);
  dff DFF_1033(CK,WX7192,WX7191);
  dff DFF_1034(CK,WX7194,WX7193);
  dff DFF_1035(CK,WX7196,WX7195);
  dff DFF_1036(CK,WX7198,WX7197);
  dff DFF_1037(CK,WX7200,WX7199);
  dff DFF_1038(CK,WX7202,WX7201);
  dff DFF_1039(CK,WX7204,WX7203);
  dff DFF_1040(CK,WX7206,WX7205);
  dff DFF_1041(CK,WX7208,WX7207);
  dff DFF_1042(CK,WX7210,WX7209);
  dff DFF_1043(CK,WX7212,WX7211);
  dff DFF_1044(CK,WX7214,WX7213);
  dff DFF_1045(CK,WX7216,WX7215);
  dff DFF_1046(CK,WX7218,WX7217);
  dff DFF_1047(CK,WX7220,WX7219);
  dff DFF_1048(CK,WX7222,WX7221);
  dff DFF_1049(CK,WX7224,WX7223);
  dff DFF_1050(CK,WX7226,WX7225);
  dff DFF_1051(CK,WX7228,WX7227);
  dff DFF_1052(CK,WX7230,WX7229);
  dff DFF_1053(CK,WX7232,WX7231);
  dff DFF_1054(CK,WX7234,WX7233);
  dff DFF_1055(CK,WX7236,WX7235);
  dff DFF_1056(CK,WX7238,WX7237);
  dff DFF_1057(CK,WX7240,WX7239);
  dff DFF_1058(CK,WX7242,WX7241);
  dff DFF_1059(CK,WX7244,WX7243);
  dff DFF_1060(CK,WX7246,WX7245);
  dff DFF_1061(CK,WX7248,WX7247);
  dff DFF_1062(CK,WX7250,WX7249);
  dff DFF_1063(CK,WX7252,WX7251);
  dff DFF_1064(CK,WX7254,WX7253);
  dff DFF_1065(CK,WX7256,WX7255);
  dff DFF_1066(CK,WX7258,WX7257);
  dff DFF_1067(CK,WX7260,WX7259);
  dff DFF_1068(CK,WX7262,WX7261);
  dff DFF_1069(CK,WX7264,WX7263);
  dff DFF_1070(CK,WX7266,WX7265);
  dff DFF_1071(CK,WX7268,WX7267);
  dff DFF_1072(CK,WX7270,WX7269);
  dff DFF_1073(CK,WX7272,WX7271);
  dff DFF_1074(CK,WX7274,WX7273);
  dff DFF_1075(CK,WX7276,WX7275);
  dff DFF_1076(CK,WX7278,WX7277);
  dff DFF_1077(CK,WX7280,WX7279);
  dff DFF_1078(CK,WX7282,WX7281);
  dff DFF_1079(CK,WX7284,WX7283);
  dff DFF_1080(CK,WX7286,WX7285);
  dff DFF_1081(CK,WX7288,WX7287);
  dff DFF_1082(CK,WX7290,WX7289);
  dff DFF_1083(CK,WX7292,WX7291);
  dff DFF_1084(CK,WX7294,WX7293);
  dff DFF_1085(CK,WX7296,WX7295);
  dff DFF_1086(CK,WX7298,WX7297);
  dff DFF_1087(CK,WX7300,WX7299);
  dff DFF_1088(CK,WX7302,WX7301);
  dff DFF_1089(CK,WX7304,WX7303);
  dff DFF_1090(CK,WX7306,WX7305);
  dff DFF_1091(CK,WX7308,WX7307);
  dff DFF_1092(CK,WX7310,WX7309);
  dff DFF_1093(CK,WX7312,WX7311);
  dff DFF_1094(CK,WX7314,WX7313);
  dff DFF_1095(CK,WX7316,WX7315);
  dff DFF_1096(CK,WX7318,WX7317);
  dff DFF_1097(CK,WX7320,WX7319);
  dff DFF_1098(CK,WX7322,WX7321);
  dff DFF_1099(CK,WX7324,WX7323);
  dff DFF_1100(CK,WX7326,WX7325);
  dff DFF_1101(CK,WX7328,WX7327);
  dff DFF_1102(CK,WX7330,WX7329);
  dff DFF_1103(CK,WX7332,WX7331);
  dff DFF_1104(CK,WX7334,WX7333);
  dff DFF_1105(CK,WX7336,WX7335);
  dff DFF_1106(CK,WX7338,WX7337);
  dff DFF_1107(CK,WX7340,WX7339);
  dff DFF_1108(CK,WX7342,WX7341);
  dff DFF_1109(CK,WX7344,WX7343);
  dff DFF_1110(CK,WX7346,WX7345);
  dff DFF_1111(CK,WX7348,WX7347);
  dff DFF_1112(CK,WX7350,WX7349);
  dff DFF_1113(CK,WX7352,WX7351);
  dff DFF_1114(CK,WX7354,WX7353);
  dff DFF_1115(CK,WX7356,WX7355);
  dff DFF_1116(CK,WX7358,WX7357);
  dff DFF_1117(CK,WX7360,WX7359);
  dff DFF_1118(CK,WX7362,WX7361);
  dff DFF_1119(CK,WX7364,WX7363);
  dff DFF_1120(CK,CRC_OUT_4_0,WX7729);
  dff DFF_1121(CK,CRC_OUT_4_1,WX7731);
  dff DFF_1122(CK,CRC_OUT_4_2,WX7733);
  dff DFF_1123(CK,CRC_OUT_4_3,WX7735);
  dff DFF_1124(CK,CRC_OUT_4_4,WX7737);
  dff DFF_1125(CK,CRC_OUT_4_5,WX7739);
  dff DFF_1126(CK,CRC_OUT_4_6,WX7741);
  dff DFF_1127(CK,CRC_OUT_4_7,WX7743);
  dff DFF_1128(CK,CRC_OUT_4_8,WX7745);
  dff DFF_1129(CK,CRC_OUT_4_9,WX7747);
  dff DFF_1130(CK,CRC_OUT_4_10,WX7749);
  dff DFF_1131(CK,CRC_OUT_4_11,WX7751);
  dff DFF_1132(CK,CRC_OUT_4_12,WX7753);
  dff DFF_1133(CK,CRC_OUT_4_13,WX7755);
  dff DFF_1134(CK,CRC_OUT_4_14,WX7757);
  dff DFF_1135(CK,CRC_OUT_4_15,WX7759);
  dff DFF_1136(CK,CRC_OUT_4_16,WX7761);
  dff DFF_1137(CK,CRC_OUT_4_17,WX7763);
  dff DFF_1138(CK,CRC_OUT_4_18,WX7765);
  dff DFF_1139(CK,CRC_OUT_4_19,WX7767);
  dff DFF_1140(CK,CRC_OUT_4_20,WX7769);
  dff DFF_1141(CK,CRC_OUT_4_21,WX7771);
  dff DFF_1142(CK,CRC_OUT_4_22,WX7773);
  dff DFF_1143(CK,CRC_OUT_4_23,WX7775);
  dff DFF_1144(CK,CRC_OUT_4_24,WX7777);
  dff DFF_1145(CK,CRC_OUT_4_25,WX7779);
  dff DFF_1146(CK,CRC_OUT_4_26,WX7781);
  dff DFF_1147(CK,CRC_OUT_4_27,WX7783);
  dff DFF_1148(CK,CRC_OUT_4_28,WX7785);
  dff DFF_1149(CK,CRC_OUT_4_29,WX7787);
  dff DFF_1150(CK,CRC_OUT_4_30,WX7789);
  dff DFF_1151(CK,CRC_OUT_4_31,WX7791);
  dff DFF_1152(CK,WX8243,WX8242);
  dff DFF_1153(CK,WX8245,WX8244);
  dff DFF_1154(CK,WX8247,WX8246);
  dff DFF_1155(CK,WX8249,WX8248);
  dff DFF_1156(CK,WX8251,WX8250);
  dff DFF_1157(CK,WX8253,WX8252);
  dff DFF_1158(CK,WX8255,WX8254);
  dff DFF_1159(CK,WX8257,WX8256);
  dff DFF_1160(CK,WX8259,WX8258);
  dff DFF_1161(CK,WX8261,WX8260);
  dff DFF_1162(CK,WX8263,WX8262);
  dff DFF_1163(CK,WX8265,WX8264);
  dff DFF_1164(CK,WX8267,WX8266);
  dff DFF_1165(CK,WX8269,WX8268);
  dff DFF_1166(CK,WX8271,WX8270);
  dff DFF_1167(CK,WX8273,WX8272);
  dff DFF_1168(CK,WX8275,WX8274);
  dff DFF_1169(CK,WX8277,WX8276);
  dff DFF_1170(CK,WX8279,WX8278);
  dff DFF_1171(CK,WX8281,WX8280);
  dff DFF_1172(CK,WX8283,WX8282);
  dff DFF_1173(CK,WX8285,WX8284);
  dff DFF_1174(CK,WX8287,WX8286);
  dff DFF_1175(CK,WX8289,WX8288);
  dff DFF_1176(CK,WX8291,WX8290);
  dff DFF_1177(CK,WX8293,WX8292);
  dff DFF_1178(CK,WX8295,WX8294);
  dff DFF_1179(CK,WX8297,WX8296);
  dff DFF_1180(CK,WX8299,WX8298);
  dff DFF_1181(CK,WX8301,WX8300);
  dff DFF_1182(CK,WX8303,WX8302);
  dff DFF_1183(CK,WX8305,WX8304);
  dff DFF_1184(CK,WX8403,WX8402);
  dff DFF_1185(CK,WX8405,WX8404);
  dff DFF_1186(CK,WX8407,WX8406);
  dff DFF_1187(CK,WX8409,WX8408);
  dff DFF_1188(CK,WX8411,WX8410);
  dff DFF_1189(CK,WX8413,WX8412);
  dff DFF_1190(CK,WX8415,WX8414);
  dff DFF_1191(CK,WX8417,WX8416);
  dff DFF_1192(CK,WX8419,WX8418);
  dff DFF_1193(CK,WX8421,WX8420);
  dff DFF_1194(CK,WX8423,WX8422);
  dff DFF_1195(CK,WX8425,WX8424);
  dff DFF_1196(CK,WX8427,WX8426);
  dff DFF_1197(CK,WX8429,WX8428);
  dff DFF_1198(CK,WX8431,WX8430);
  dff DFF_1199(CK,WX8433,WX8432);
  dff DFF_1200(CK,WX8435,WX8434);
  dff DFF_1201(CK,WX8437,WX8436);
  dff DFF_1202(CK,WX8439,WX8438);
  dff DFF_1203(CK,WX8441,WX8440);
  dff DFF_1204(CK,WX8443,WX8442);
  dff DFF_1205(CK,WX8445,WX8444);
  dff DFF_1206(CK,WX8447,WX8446);
  dff DFF_1207(CK,WX8449,WX8448);
  dff DFF_1208(CK,WX8451,WX8450);
  dff DFF_1209(CK,WX8453,WX8452);
  dff DFF_1210(CK,WX8455,WX8454);
  dff DFF_1211(CK,WX8457,WX8456);
  dff DFF_1212(CK,WX8459,WX8458);
  dff DFF_1213(CK,WX8461,WX8460);
  dff DFF_1214(CK,WX8463,WX8462);
  dff DFF_1215(CK,WX8465,WX8464);
  dff DFF_1216(CK,WX8467,WX8466);
  dff DFF_1217(CK,WX8469,WX8468);
  dff DFF_1218(CK,WX8471,WX8470);
  dff DFF_1219(CK,WX8473,WX8472);
  dff DFF_1220(CK,WX8475,WX8474);
  dff DFF_1221(CK,WX8477,WX8476);
  dff DFF_1222(CK,WX8479,WX8478);
  dff DFF_1223(CK,WX8481,WX8480);
  dff DFF_1224(CK,WX8483,WX8482);
  dff DFF_1225(CK,WX8485,WX8484);
  dff DFF_1226(CK,WX8487,WX8486);
  dff DFF_1227(CK,WX8489,WX8488);
  dff DFF_1228(CK,WX8491,WX8490);
  dff DFF_1229(CK,WX8493,WX8492);
  dff DFF_1230(CK,WX8495,WX8494);
  dff DFF_1231(CK,WX8497,WX8496);
  dff DFF_1232(CK,WX8499,WX8498);
  dff DFF_1233(CK,WX8501,WX8500);
  dff DFF_1234(CK,WX8503,WX8502);
  dff DFF_1235(CK,WX8505,WX8504);
  dff DFF_1236(CK,WX8507,WX8506);
  dff DFF_1237(CK,WX8509,WX8508);
  dff DFF_1238(CK,WX8511,WX8510);
  dff DFF_1239(CK,WX8513,WX8512);
  dff DFF_1240(CK,WX8515,WX8514);
  dff DFF_1241(CK,WX8517,WX8516);
  dff DFF_1242(CK,WX8519,WX8518);
  dff DFF_1243(CK,WX8521,WX8520);
  dff DFF_1244(CK,WX8523,WX8522);
  dff DFF_1245(CK,WX8525,WX8524);
  dff DFF_1246(CK,WX8527,WX8526);
  dff DFF_1247(CK,WX8529,WX8528);
  dff DFF_1248(CK,WX8531,WX8530);
  dff DFF_1249(CK,WX8533,WX8532);
  dff DFF_1250(CK,WX8535,WX8534);
  dff DFF_1251(CK,WX8537,WX8536);
  dff DFF_1252(CK,WX8539,WX8538);
  dff DFF_1253(CK,WX8541,WX8540);
  dff DFF_1254(CK,WX8543,WX8542);
  dff DFF_1255(CK,WX8545,WX8544);
  dff DFF_1256(CK,WX8547,WX8546);
  dff DFF_1257(CK,WX8549,WX8548);
  dff DFF_1258(CK,WX8551,WX8550);
  dff DFF_1259(CK,WX8553,WX8552);
  dff DFF_1260(CK,WX8555,WX8554);
  dff DFF_1261(CK,WX8557,WX8556);
  dff DFF_1262(CK,WX8559,WX8558);
  dff DFF_1263(CK,WX8561,WX8560);
  dff DFF_1264(CK,WX8563,WX8562);
  dff DFF_1265(CK,WX8565,WX8564);
  dff DFF_1266(CK,WX8567,WX8566);
  dff DFF_1267(CK,WX8569,WX8568);
  dff DFF_1268(CK,WX8571,WX8570);
  dff DFF_1269(CK,WX8573,WX8572);
  dff DFF_1270(CK,WX8575,WX8574);
  dff DFF_1271(CK,WX8577,WX8576);
  dff DFF_1272(CK,WX8579,WX8578);
  dff DFF_1273(CK,WX8581,WX8580);
  dff DFF_1274(CK,WX8583,WX8582);
  dff DFF_1275(CK,WX8585,WX8584);
  dff DFF_1276(CK,WX8587,WX8586);
  dff DFF_1277(CK,WX8589,WX8588);
  dff DFF_1278(CK,WX8591,WX8590);
  dff DFF_1279(CK,WX8593,WX8592);
  dff DFF_1280(CK,WX8595,WX8594);
  dff DFF_1281(CK,WX8597,WX8596);
  dff DFF_1282(CK,WX8599,WX8598);
  dff DFF_1283(CK,WX8601,WX8600);
  dff DFF_1284(CK,WX8603,WX8602);
  dff DFF_1285(CK,WX8605,WX8604);
  dff DFF_1286(CK,WX8607,WX8606);
  dff DFF_1287(CK,WX8609,WX8608);
  dff DFF_1288(CK,WX8611,WX8610);
  dff DFF_1289(CK,WX8613,WX8612);
  dff DFF_1290(CK,WX8615,WX8614);
  dff DFF_1291(CK,WX8617,WX8616);
  dff DFF_1292(CK,WX8619,WX8618);
  dff DFF_1293(CK,WX8621,WX8620);
  dff DFF_1294(CK,WX8623,WX8622);
  dff DFF_1295(CK,WX8625,WX8624);
  dff DFF_1296(CK,WX8627,WX8626);
  dff DFF_1297(CK,WX8629,WX8628);
  dff DFF_1298(CK,WX8631,WX8630);
  dff DFF_1299(CK,WX8633,WX8632);
  dff DFF_1300(CK,WX8635,WX8634);
  dff DFF_1301(CK,WX8637,WX8636);
  dff DFF_1302(CK,WX8639,WX8638);
  dff DFF_1303(CK,WX8641,WX8640);
  dff DFF_1304(CK,WX8643,WX8642);
  dff DFF_1305(CK,WX8645,WX8644);
  dff DFF_1306(CK,WX8647,WX8646);
  dff DFF_1307(CK,WX8649,WX8648);
  dff DFF_1308(CK,WX8651,WX8650);
  dff DFF_1309(CK,WX8653,WX8652);
  dff DFF_1310(CK,WX8655,WX8654);
  dff DFF_1311(CK,WX8657,WX8656);
  dff DFF_1312(CK,CRC_OUT_3_0,WX9022);
  dff DFF_1313(CK,CRC_OUT_3_1,WX9024);
  dff DFF_1314(CK,CRC_OUT_3_2,WX9026);
  dff DFF_1315(CK,CRC_OUT_3_3,WX9028);
  dff DFF_1316(CK,CRC_OUT_3_4,WX9030);
  dff DFF_1317(CK,CRC_OUT_3_5,WX9032);
  dff DFF_1318(CK,CRC_OUT_3_6,WX9034);
  dff DFF_1319(CK,CRC_OUT_3_7,WX9036);
  dff DFF_1320(CK,CRC_OUT_3_8,WX9038);
  dff DFF_1321(CK,CRC_OUT_3_9,WX9040);
  dff DFF_1322(CK,CRC_OUT_3_10,WX9042);
  dff DFF_1323(CK,CRC_OUT_3_11,WX9044);
  dff DFF_1324(CK,CRC_OUT_3_12,WX9046);
  dff DFF_1325(CK,CRC_OUT_3_13,WX9048);
  dff DFF_1326(CK,CRC_OUT_3_14,WX9050);
  dff DFF_1327(CK,CRC_OUT_3_15,WX9052);
  dff DFF_1328(CK,CRC_OUT_3_16,WX9054);
  dff DFF_1329(CK,CRC_OUT_3_17,WX9056);
  dff DFF_1330(CK,CRC_OUT_3_18,WX9058);
  dff DFF_1331(CK,CRC_OUT_3_19,WX9060);
  dff DFF_1332(CK,CRC_OUT_3_20,WX9062);
  dff DFF_1333(CK,CRC_OUT_3_21,WX9064);
  dff DFF_1334(CK,CRC_OUT_3_22,WX9066);
  dff DFF_1335(CK,CRC_OUT_3_23,WX9068);
  dff DFF_1336(CK,CRC_OUT_3_24,WX9070);
  dff DFF_1337(CK,CRC_OUT_3_25,WX9072);
  dff DFF_1338(CK,CRC_OUT_3_26,WX9074);
  dff DFF_1339(CK,CRC_OUT_3_27,WX9076);
  dff DFF_1340(CK,CRC_OUT_3_28,WX9078);
  dff DFF_1341(CK,CRC_OUT_3_29,WX9080);
  dff DFF_1342(CK,CRC_OUT_3_30,WX9082);
  dff DFF_1343(CK,CRC_OUT_3_31,WX9084);
  dff DFF_1344(CK,WX9536,WX9535);
  dff DFF_1345(CK,WX9538,WX9537);
  dff DFF_1346(CK,WX9540,WX9539);
  dff DFF_1347(CK,WX9542,WX9541);
  dff DFF_1348(CK,WX9544,WX9543);
  dff DFF_1349(CK,WX9546,WX9545);
  dff DFF_1350(CK,WX9548,WX9547);
  dff DFF_1351(CK,WX9550,WX9549);
  dff DFF_1352(CK,WX9552,WX9551);
  dff DFF_1353(CK,WX9554,WX9553);
  dff DFF_1354(CK,WX9556,WX9555);
  dff DFF_1355(CK,WX9558,WX9557);
  dff DFF_1356(CK,WX9560,WX9559);
  dff DFF_1357(CK,WX9562,WX9561);
  dff DFF_1358(CK,WX9564,WX9563);
  dff DFF_1359(CK,WX9566,WX9565);
  dff DFF_1360(CK,WX9568,WX9567);
  dff DFF_1361(CK,WX9570,WX9569);
  dff DFF_1362(CK,WX9572,WX9571);
  dff DFF_1363(CK,WX9574,WX9573);
  dff DFF_1364(CK,WX9576,WX9575);
  dff DFF_1365(CK,WX9578,WX9577);
  dff DFF_1366(CK,WX9580,WX9579);
  dff DFF_1367(CK,WX9582,WX9581);
  dff DFF_1368(CK,WX9584,WX9583);
  dff DFF_1369(CK,WX9586,WX9585);
  dff DFF_1370(CK,WX9588,WX9587);
  dff DFF_1371(CK,WX9590,WX9589);
  dff DFF_1372(CK,WX9592,WX9591);
  dff DFF_1373(CK,WX9594,WX9593);
  dff DFF_1374(CK,WX9596,WX9595);
  dff DFF_1375(CK,WX9598,WX9597);
  dff DFF_1376(CK,WX9696,WX9695);
  dff DFF_1377(CK,WX9698,WX9697);
  dff DFF_1378(CK,WX9700,WX9699);
  dff DFF_1379(CK,WX9702,WX9701);
  dff DFF_1380(CK,WX9704,WX9703);
  dff DFF_1381(CK,WX9706,WX9705);
  dff DFF_1382(CK,WX9708,WX9707);
  dff DFF_1383(CK,WX9710,WX9709);
  dff DFF_1384(CK,WX9712,WX9711);
  dff DFF_1385(CK,WX9714,WX9713);
  dff DFF_1386(CK,WX9716,WX9715);
  dff DFF_1387(CK,WX9718,WX9717);
  dff DFF_1388(CK,WX9720,WX9719);
  dff DFF_1389(CK,WX9722,WX9721);
  dff DFF_1390(CK,WX9724,WX9723);
  dff DFF_1391(CK,WX9726,WX9725);
  dff DFF_1392(CK,WX9728,WX9727);
  dff DFF_1393(CK,WX9730,WX9729);
  dff DFF_1394(CK,WX9732,WX9731);
  dff DFF_1395(CK,WX9734,WX9733);
  dff DFF_1396(CK,WX9736,WX9735);
  dff DFF_1397(CK,WX9738,WX9737);
  dff DFF_1398(CK,WX9740,WX9739);
  dff DFF_1399(CK,WX9742,WX9741);
  dff DFF_1400(CK,WX9744,WX9743);
  dff DFF_1401(CK,WX9746,WX9745);
  dff DFF_1402(CK,WX9748,WX9747);
  dff DFF_1403(CK,WX9750,WX9749);
  dff DFF_1404(CK,WX9752,WX9751);
  dff DFF_1405(CK,WX9754,WX9753);
  dff DFF_1406(CK,WX9756,WX9755);
  dff DFF_1407(CK,WX9758,WX9757);
  dff DFF_1408(CK,WX9760,WX9759);
  dff DFF_1409(CK,WX9762,WX9761);
  dff DFF_1410(CK,WX9764,WX9763);
  dff DFF_1411(CK,WX9766,WX9765);
  dff DFF_1412(CK,WX9768,WX9767);
  dff DFF_1413(CK,WX9770,WX9769);
  dff DFF_1414(CK,WX9772,WX9771);
  dff DFF_1415(CK,WX9774,WX9773);
  dff DFF_1416(CK,WX9776,WX9775);
  dff DFF_1417(CK,WX9778,WX9777);
  dff DFF_1418(CK,WX9780,WX9779);
  dff DFF_1419(CK,WX9782,WX9781);
  dff DFF_1420(CK,WX9784,WX9783);
  dff DFF_1421(CK,WX9786,WX9785);
  dff DFF_1422(CK,WX9788,WX9787);
  dff DFF_1423(CK,WX9790,WX9789);
  dff DFF_1424(CK,WX9792,WX9791);
  dff DFF_1425(CK,WX9794,WX9793);
  dff DFF_1426(CK,WX9796,WX9795);
  dff DFF_1427(CK,WX9798,WX9797);
  dff DFF_1428(CK,WX9800,WX9799);
  dff DFF_1429(CK,WX9802,WX9801);
  dff DFF_1430(CK,WX9804,WX9803);
  dff DFF_1431(CK,WX9806,WX9805);
  dff DFF_1432(CK,WX9808,WX9807);
  dff DFF_1433(CK,WX9810,WX9809);
  dff DFF_1434(CK,WX9812,WX9811);
  dff DFF_1435(CK,WX9814,WX9813);
  dff DFF_1436(CK,WX9816,WX9815);
  dff DFF_1437(CK,WX9818,WX9817);
  dff DFF_1438(CK,WX9820,WX9819);
  dff DFF_1439(CK,WX9822,WX9821);
  dff DFF_1440(CK,WX9824,WX9823);
  dff DFF_1441(CK,WX9826,WX9825);
  dff DFF_1442(CK,WX9828,WX9827);
  dff DFF_1443(CK,WX9830,WX9829);
  dff DFF_1444(CK,WX9832,WX9831);
  dff DFF_1445(CK,WX9834,WX9833);
  dff DFF_1446(CK,WX9836,WX9835);
  dff DFF_1447(CK,WX9838,WX9837);
  dff DFF_1448(CK,WX9840,WX9839);
  dff DFF_1449(CK,WX9842,WX9841);
  dff DFF_1450(CK,WX9844,WX9843);
  dff DFF_1451(CK,WX9846,WX9845);
  dff DFF_1452(CK,WX9848,WX9847);
  dff DFF_1453(CK,WX9850,WX9849);
  dff DFF_1454(CK,WX9852,WX9851);
  dff DFF_1455(CK,WX9854,WX9853);
  dff DFF_1456(CK,WX9856,WX9855);
  dff DFF_1457(CK,WX9858,WX9857);
  dff DFF_1458(CK,WX9860,WX9859);
  dff DFF_1459(CK,WX9862,WX9861);
  dff DFF_1460(CK,WX9864,WX9863);
  dff DFF_1461(CK,WX9866,WX9865);
  dff DFF_1462(CK,WX9868,WX9867);
  dff DFF_1463(CK,WX9870,WX9869);
  dff DFF_1464(CK,WX9872,WX9871);
  dff DFF_1465(CK,WX9874,WX9873);
  dff DFF_1466(CK,WX9876,WX9875);
  dff DFF_1467(CK,WX9878,WX9877);
  dff DFF_1468(CK,WX9880,WX9879);
  dff DFF_1469(CK,WX9882,WX9881);
  dff DFF_1470(CK,WX9884,WX9883);
  dff DFF_1471(CK,WX9886,WX9885);
  dff DFF_1472(CK,WX9888,WX9887);
  dff DFF_1473(CK,WX9890,WX9889);
  dff DFF_1474(CK,WX9892,WX9891);
  dff DFF_1475(CK,WX9894,WX9893);
  dff DFF_1476(CK,WX9896,WX9895);
  dff DFF_1477(CK,WX9898,WX9897);
  dff DFF_1478(CK,WX9900,WX9899);
  dff DFF_1479(CK,WX9902,WX9901);
  dff DFF_1480(CK,WX9904,WX9903);
  dff DFF_1481(CK,WX9906,WX9905);
  dff DFF_1482(CK,WX9908,WX9907);
  dff DFF_1483(CK,WX9910,WX9909);
  dff DFF_1484(CK,WX9912,WX9911);
  dff DFF_1485(CK,WX9914,WX9913);
  dff DFF_1486(CK,WX9916,WX9915);
  dff DFF_1487(CK,WX9918,WX9917);
  dff DFF_1488(CK,WX9920,WX9919);
  dff DFF_1489(CK,WX9922,WX9921);
  dff DFF_1490(CK,WX9924,WX9923);
  dff DFF_1491(CK,WX9926,WX9925);
  dff DFF_1492(CK,WX9928,WX9927);
  dff DFF_1493(CK,WX9930,WX9929);
  dff DFF_1494(CK,WX9932,WX9931);
  dff DFF_1495(CK,WX9934,WX9933);
  dff DFF_1496(CK,WX9936,WX9935);
  dff DFF_1497(CK,WX9938,WX9937);
  dff DFF_1498(CK,WX9940,WX9939);
  dff DFF_1499(CK,WX9942,WX9941);
  dff DFF_1500(CK,WX9944,WX9943);
  dff DFF_1501(CK,WX9946,WX9945);
  dff DFF_1502(CK,WX9948,WX9947);
  dff DFF_1503(CK,WX9950,WX9949);
  dff DFF_1504(CK,CRC_OUT_2_0,WX10315);
  dff DFF_1505(CK,CRC_OUT_2_1,WX10317);
  dff DFF_1506(CK,CRC_OUT_2_2,WX10319);
  dff DFF_1507(CK,CRC_OUT_2_3,WX10321);
  dff DFF_1508(CK,CRC_OUT_2_4,WX10323);
  dff DFF_1509(CK,CRC_OUT_2_5,WX10325);
  dff DFF_1510(CK,CRC_OUT_2_6,WX10327);
  dff DFF_1511(CK,CRC_OUT_2_7,WX10329);
  dff DFF_1512(CK,CRC_OUT_2_8,WX10331);
  dff DFF_1513(CK,CRC_OUT_2_9,WX10333);
  dff DFF_1514(CK,CRC_OUT_2_10,WX10335);
  dff DFF_1515(CK,CRC_OUT_2_11,WX10337);
  dff DFF_1516(CK,CRC_OUT_2_12,WX10339);
  dff DFF_1517(CK,CRC_OUT_2_13,WX10341);
  dff DFF_1518(CK,CRC_OUT_2_14,WX10343);
  dff DFF_1519(CK,CRC_OUT_2_15,WX10345);
  dff DFF_1520(CK,CRC_OUT_2_16,WX10347);
  dff DFF_1521(CK,CRC_OUT_2_17,WX10349);
  dff DFF_1522(CK,CRC_OUT_2_18,WX10351);
  dff DFF_1523(CK,CRC_OUT_2_19,WX10353);
  dff DFF_1524(CK,CRC_OUT_2_20,WX10355);
  dff DFF_1525(CK,CRC_OUT_2_21,WX10357);
  dff DFF_1526(CK,CRC_OUT_2_22,WX10359);
  dff DFF_1527(CK,CRC_OUT_2_23,WX10361);
  dff DFF_1528(CK,CRC_OUT_2_24,WX10363);
  dff DFF_1529(CK,CRC_OUT_2_25,WX10365);
  dff DFF_1530(CK,CRC_OUT_2_26,WX10367);
  dff DFF_1531(CK,CRC_OUT_2_27,WX10369);
  dff DFF_1532(CK,CRC_OUT_2_28,WX10371);
  dff DFF_1533(CK,CRC_OUT_2_29,WX10373);
  dff DFF_1534(CK,CRC_OUT_2_30,WX10375);
  dff DFF_1535(CK,CRC_OUT_2_31,WX10377);
  dff DFF_1536(CK,WX10829,WX10828);
  dff DFF_1537(CK,WX10831,WX10830);
  dff DFF_1538(CK,WX10833,WX10832);
  dff DFF_1539(CK,WX10835,WX10834);
  dff DFF_1540(CK,WX10837,WX10836);
  dff DFF_1541(CK,WX10839,WX10838);
  dff DFF_1542(CK,WX10841,WX10840);
  dff DFF_1543(CK,WX10843,WX10842);
  dff DFF_1544(CK,WX10845,WX10844);
  dff DFF_1545(CK,WX10847,WX10846);
  dff DFF_1546(CK,WX10849,WX10848);
  dff DFF_1547(CK,WX10851,WX10850);
  dff DFF_1548(CK,WX10853,WX10852);
  dff DFF_1549(CK,WX10855,WX10854);
  dff DFF_1550(CK,WX10857,WX10856);
  dff DFF_1551(CK,WX10859,WX10858);
  dff DFF_1552(CK,WX10861,WX10860);
  dff DFF_1553(CK,WX10863,WX10862);
  dff DFF_1554(CK,WX10865,WX10864);
  dff DFF_1555(CK,WX10867,WX10866);
  dff DFF_1556(CK,WX10869,WX10868);
  dff DFF_1557(CK,WX10871,WX10870);
  dff DFF_1558(CK,WX10873,WX10872);
  dff DFF_1559(CK,WX10875,WX10874);
  dff DFF_1560(CK,WX10877,WX10876);
  dff DFF_1561(CK,WX10879,WX10878);
  dff DFF_1562(CK,WX10881,WX10880);
  dff DFF_1563(CK,WX10883,WX10882);
  dff DFF_1564(CK,WX10885,WX10884);
  dff DFF_1565(CK,WX10887,WX10886);
  dff DFF_1566(CK,WX10889,WX10888);
  dff DFF_1567(CK,WX10891,WX10890);
  dff DFF_1568(CK,WX10989,WX10988);
  dff DFF_1569(CK,WX10991,WX10990);
  dff DFF_1570(CK,WX10993,WX10992);
  dff DFF_1571(CK,WX10995,WX10994);
  dff DFF_1572(CK,WX10997,WX10996);
  dff DFF_1573(CK,WX10999,WX10998);
  dff DFF_1574(CK,WX11001,WX11000);
  dff DFF_1575(CK,WX11003,WX11002);
  dff DFF_1576(CK,WX11005,WX11004);
  dff DFF_1577(CK,WX11007,WX11006);
  dff DFF_1578(CK,WX11009,WX11008);
  dff DFF_1579(CK,WX11011,WX11010);
  dff DFF_1580(CK,WX11013,WX11012);
  dff DFF_1581(CK,WX11015,WX11014);
  dff DFF_1582(CK,WX11017,WX11016);
  dff DFF_1583(CK,WX11019,WX11018);
  dff DFF_1584(CK,WX11021,WX11020);
  dff DFF_1585(CK,WX11023,WX11022);
  dff DFF_1586(CK,WX11025,WX11024);
  dff DFF_1587(CK,WX11027,WX11026);
  dff DFF_1588(CK,WX11029,WX11028);
  dff DFF_1589(CK,WX11031,WX11030);
  dff DFF_1590(CK,WX11033,WX11032);
  dff DFF_1591(CK,WX11035,WX11034);
  dff DFF_1592(CK,WX11037,WX11036);
  dff DFF_1593(CK,WX11039,WX11038);
  dff DFF_1594(CK,WX11041,WX11040);
  dff DFF_1595(CK,WX11043,WX11042);
  dff DFF_1596(CK,WX11045,WX11044);
  dff DFF_1597(CK,WX11047,WX11046);
  dff DFF_1598(CK,WX11049,WX11048);
  dff DFF_1599(CK,WX11051,WX11050);
  dff DFF_1600(CK,WX11053,WX11052);
  dff DFF_1601(CK,WX11055,WX11054);
  dff DFF_1602(CK,WX11057,WX11056);
  dff DFF_1603(CK,WX11059,WX11058);
  dff DFF_1604(CK,WX11061,WX11060);
  dff DFF_1605(CK,WX11063,WX11062);
  dff DFF_1606(CK,WX11065,WX11064);
  dff DFF_1607(CK,WX11067,WX11066);
  dff DFF_1608(CK,WX11069,WX11068);
  dff DFF_1609(CK,WX11071,WX11070);
  dff DFF_1610(CK,WX11073,WX11072);
  dff DFF_1611(CK,WX11075,WX11074);
  dff DFF_1612(CK,WX11077,WX11076);
  dff DFF_1613(CK,WX11079,WX11078);
  dff DFF_1614(CK,WX11081,WX11080);
  dff DFF_1615(CK,WX11083,WX11082);
  dff DFF_1616(CK,WX11085,WX11084);
  dff DFF_1617(CK,WX11087,WX11086);
  dff DFF_1618(CK,WX11089,WX11088);
  dff DFF_1619(CK,WX11091,WX11090);
  dff DFF_1620(CK,WX11093,WX11092);
  dff DFF_1621(CK,WX11095,WX11094);
  dff DFF_1622(CK,WX11097,WX11096);
  dff DFF_1623(CK,WX11099,WX11098);
  dff DFF_1624(CK,WX11101,WX11100);
  dff DFF_1625(CK,WX11103,WX11102);
  dff DFF_1626(CK,WX11105,WX11104);
  dff DFF_1627(CK,WX11107,WX11106);
  dff DFF_1628(CK,WX11109,WX11108);
  dff DFF_1629(CK,WX11111,WX11110);
  dff DFF_1630(CK,WX11113,WX11112);
  dff DFF_1631(CK,WX11115,WX11114);
  dff DFF_1632(CK,WX11117,WX11116);
  dff DFF_1633(CK,WX11119,WX11118);
  dff DFF_1634(CK,WX11121,WX11120);
  dff DFF_1635(CK,WX11123,WX11122);
  dff DFF_1636(CK,WX11125,WX11124);
  dff DFF_1637(CK,WX11127,WX11126);
  dff DFF_1638(CK,WX11129,WX11128);
  dff DFF_1639(CK,WX11131,WX11130);
  dff DFF_1640(CK,WX11133,WX11132);
  dff DFF_1641(CK,WX11135,WX11134);
  dff DFF_1642(CK,WX11137,WX11136);
  dff DFF_1643(CK,WX11139,WX11138);
  dff DFF_1644(CK,WX11141,WX11140);
  dff DFF_1645(CK,WX11143,WX11142);
  dff DFF_1646(CK,WX11145,WX11144);
  dff DFF_1647(CK,WX11147,WX11146);
  dff DFF_1648(CK,WX11149,WX11148);
  dff DFF_1649(CK,WX11151,WX11150);
  dff DFF_1650(CK,WX11153,WX11152);
  dff DFF_1651(CK,WX11155,WX11154);
  dff DFF_1652(CK,WX11157,WX11156);
  dff DFF_1653(CK,WX11159,WX11158);
  dff DFF_1654(CK,WX11161,WX11160);
  dff DFF_1655(CK,WX11163,WX11162);
  dff DFF_1656(CK,WX11165,WX11164);
  dff DFF_1657(CK,WX11167,WX11166);
  dff DFF_1658(CK,WX11169,WX11168);
  dff DFF_1659(CK,WX11171,WX11170);
  dff DFF_1660(CK,WX11173,WX11172);
  dff DFF_1661(CK,WX11175,WX11174);
  dff DFF_1662(CK,WX11177,WX11176);
  dff DFF_1663(CK,WX11179,WX11178);
  dff DFF_1664(CK,WX11181,WX11180);
  dff DFF_1665(CK,WX11183,WX11182);
  dff DFF_1666(CK,WX11185,WX11184);
  dff DFF_1667(CK,WX11187,WX11186);
  dff DFF_1668(CK,WX11189,WX11188);
  dff DFF_1669(CK,WX11191,WX11190);
  dff DFF_1670(CK,WX11193,WX11192);
  dff DFF_1671(CK,WX11195,WX11194);
  dff DFF_1672(CK,WX11197,WX11196);
  dff DFF_1673(CK,WX11199,WX11198);
  dff DFF_1674(CK,WX11201,WX11200);
  dff DFF_1675(CK,WX11203,WX11202);
  dff DFF_1676(CK,WX11205,WX11204);
  dff DFF_1677(CK,WX11207,WX11206);
  dff DFF_1678(CK,WX11209,WX11208);
  dff DFF_1679(CK,WX11211,WX11210);
  dff DFF_1680(CK,WX11213,WX11212);
  dff DFF_1681(CK,WX11215,WX11214);
  dff DFF_1682(CK,WX11217,WX11216);
  dff DFF_1683(CK,WX11219,WX11218);
  dff DFF_1684(CK,WX11221,WX11220);
  dff DFF_1685(CK,WX11223,WX11222);
  dff DFF_1686(CK,WX11225,WX11224);
  dff DFF_1687(CK,WX11227,WX11226);
  dff DFF_1688(CK,WX11229,WX11228);
  dff DFF_1689(CK,WX11231,WX11230);
  dff DFF_1690(CK,WX11233,WX11232);
  dff DFF_1691(CK,WX11235,WX11234);
  dff DFF_1692(CK,WX11237,WX11236);
  dff DFF_1693(CK,WX11239,WX11238);
  dff DFF_1694(CK,WX11241,WX11240);
  dff DFF_1695(CK,WX11243,WX11242);
  dff DFF_1696(CK,CRC_OUT_1_0,WX11608);
  dff DFF_1697(CK,CRC_OUT_1_1,WX11610);
  dff DFF_1698(CK,CRC_OUT_1_2,WX11612);
  dff DFF_1699(CK,CRC_OUT_1_3,WX11614);
  dff DFF_1700(CK,CRC_OUT_1_4,WX11616);
  dff DFF_1701(CK,CRC_OUT_1_5,WX11618);
  dff DFF_1702(CK,CRC_OUT_1_6,WX11620);
  dff DFF_1703(CK,CRC_OUT_1_7,WX11622);
  dff DFF_1704(CK,CRC_OUT_1_8,WX11624);
  dff DFF_1705(CK,CRC_OUT_1_9,WX11626);
  dff DFF_1706(CK,CRC_OUT_1_10,WX11628);
  dff DFF_1707(CK,CRC_OUT_1_11,WX11630);
  dff DFF_1708(CK,CRC_OUT_1_12,WX11632);
  dff DFF_1709(CK,CRC_OUT_1_13,WX11634);
  dff DFF_1710(CK,CRC_OUT_1_14,WX11636);
  dff DFF_1711(CK,CRC_OUT_1_15,WX11638);
  dff DFF_1712(CK,CRC_OUT_1_16,WX11640);
  dff DFF_1713(CK,CRC_OUT_1_17,WX11642);
  dff DFF_1714(CK,CRC_OUT_1_18,WX11644);
  dff DFF_1715(CK,CRC_OUT_1_19,WX11646);
  dff DFF_1716(CK,CRC_OUT_1_20,WX11648);
  dff DFF_1717(CK,CRC_OUT_1_21,WX11650);
  dff DFF_1718(CK,CRC_OUT_1_22,WX11652);
  dff DFF_1719(CK,CRC_OUT_1_23,WX11654);
  dff DFF_1720(CK,CRC_OUT_1_24,WX11656);
  dff DFF_1721(CK,CRC_OUT_1_25,WX11658);
  dff DFF_1722(CK,CRC_OUT_1_26,WX11660);
  dff DFF_1723(CK,CRC_OUT_1_27,WX11662);
  dff DFF_1724(CK,CRC_OUT_1_28,WX11664);
  dff DFF_1725(CK,CRC_OUT_1_29,WX11666);
  dff DFF_1726(CK,CRC_OUT_1_30,WX11668);
  dff DFF_1727(CK,CRC_OUT_1_31,WX11670);
  not NOT_0(WX37,WX1003);
  not NOT_1(WX41,WX1004);
  not NOT_2(WX45,WX1004);
  not NOT_3(WX47,WX38);
  not NOT_4(WX48,WX47);
  not NOT_5(WX51,WX1003);
  not NOT_6(WX55,WX1004);
  not NOT_7(WX59,WX1004);
  not NOT_8(WX61,WX52);
  not NOT_9(WX62,WX61);
  not NOT_10(WX65,WX1003);
  not NOT_11(WX69,WX1004);
  not NOT_12(WX73,WX1004);
  not NOT_13(WX75,WX66);
  not NOT_14(WX76,WX75);
  not NOT_15(WX79,WX1003);
  not NOT_16(WX83,WX1004);
  not NOT_17(WX87,WX1004);
  not NOT_18(WX89,WX80);
  not NOT_19(WX90,WX89);
  not NOT_20(WX93,WX1003);
  not NOT_21(WX97,WX1004);
  not NOT_22(WX101,WX1004);
  not NOT_23(WX103,WX94);
  not NOT_24(WX104,WX103);
  not NOT_25(WX107,WX1003);
  not NOT_26(WX111,WX1004);
  not NOT_27(WX115,WX1004);
  not NOT_28(WX117,WX108);
  not NOT_29(WX118,WX117);
  not NOT_30(WX121,WX1003);
  not NOT_31(WX125,WX1004);
  not NOT_32(WX129,WX1004);
  not NOT_33(WX131,WX122);
  not NOT_34(WX132,WX131);
  not NOT_35(WX135,WX1003);
  not NOT_36(WX139,WX1004);
  not NOT_37(WX143,WX1004);
  not NOT_38(WX145,WX136);
  not NOT_39(WX146,WX145);
  not NOT_40(WX149,WX1003);
  not NOT_41(WX153,WX1004);
  not NOT_42(WX157,WX1004);
  not NOT_43(WX159,WX150);
  not NOT_44(WX160,WX159);
  not NOT_45(WX163,WX1003);
  not NOT_46(WX167,WX1004);
  not NOT_47(WX171,WX1004);
  not NOT_48(WX173,WX164);
  not NOT_49(WX174,WX173);
  not NOT_50(WX177,WX1003);
  not NOT_51(WX181,WX1004);
  not NOT_52(WX185,WX1004);
  not NOT_53(WX187,WX178);
  not NOT_54(WX188,WX187);
  not NOT_55(WX191,WX1003);
  not NOT_56(WX195,WX1004);
  not NOT_57(WX199,WX1004);
  not NOT_58(WX201,WX192);
  not NOT_59(WX202,WX201);
  not NOT_60(WX205,WX1003);
  not NOT_61(WX209,WX1004);
  not NOT_62(WX213,WX1004);
  not NOT_63(WX215,WX206);
  not NOT_64(WX216,WX215);
  not NOT_65(WX219,WX1003);
  not NOT_66(WX223,WX1004);
  not NOT_67(WX227,WX1004);
  not NOT_68(WX229,WX220);
  not NOT_69(WX230,WX229);
  not NOT_70(WX233,WX1003);
  not NOT_71(WX237,WX1004);
  not NOT_72(WX241,WX1004);
  not NOT_73(WX243,WX234);
  not NOT_74(WX244,WX243);
  not NOT_75(WX247,WX1003);
  not NOT_76(WX251,WX1004);
  not NOT_77(WX255,WX1004);
  not NOT_78(WX257,WX248);
  not NOT_79(WX258,WX257);
  not NOT_80(WX261,WX1003);
  not NOT_81(WX265,WX1004);
  not NOT_82(WX269,WX1004);
  not NOT_83(WX271,WX262);
  not NOT_84(WX272,WX271);
  not NOT_85(WX275,WX1003);
  not NOT_86(WX279,WX1004);
  not NOT_87(WX283,WX1004);
  not NOT_88(WX285,WX276);
  not NOT_89(WX286,WX285);
  not NOT_90(WX289,WX1003);
  not NOT_91(WX293,WX1004);
  not NOT_92(WX297,WX1004);
  not NOT_93(WX299,WX290);
  not NOT_94(WX300,WX299);
  not NOT_95(WX303,WX1003);
  not NOT_96(WX307,WX1004);
  not NOT_97(WX311,WX1004);
  not NOT_98(WX313,WX304);
  not NOT_99(WX314,WX313);
  not NOT_100(WX317,WX1003);
  not NOT_101(WX321,WX1004);
  not NOT_102(WX325,WX1004);
  not NOT_103(WX327,WX318);
  not NOT_104(WX328,WX327);
  not NOT_105(WX331,WX1003);
  not NOT_106(WX335,WX1004);
  not NOT_107(WX339,WX1004);
  not NOT_108(WX341,WX332);
  not NOT_109(WX342,WX341);
  not NOT_110(WX345,WX1003);
  not NOT_111(WX349,WX1004);
  not NOT_112(WX353,WX1004);
  not NOT_113(WX355,WX346);
  not NOT_114(WX356,WX355);
  not NOT_115(WX359,WX1003);
  not NOT_116(WX363,WX1004);
  not NOT_117(WX367,WX1004);
  not NOT_118(WX369,WX360);
  not NOT_119(WX370,WX369);
  not NOT_120(WX373,WX1003);
  not NOT_121(WX377,WX1004);
  not NOT_122(WX381,WX1004);
  not NOT_123(WX383,WX374);
  not NOT_124(WX384,WX383);
  not NOT_125(WX387,WX1003);
  not NOT_126(WX391,WX1004);
  not NOT_127(WX395,WX1004);
  not NOT_128(WX397,WX388);
  not NOT_129(WX398,WX397);
  not NOT_130(WX401,WX1003);
  not NOT_131(WX405,WX1004);
  not NOT_132(WX409,WX1004);
  not NOT_133(WX411,WX402);
  not NOT_134(WX412,WX411);
  not NOT_135(WX415,WX1003);
  not NOT_136(WX419,WX1004);
  not NOT_137(WX423,WX1004);
  not NOT_138(WX425,WX416);
  not NOT_139(WX426,WX425);
  not NOT_140(WX429,WX1003);
  not NOT_141(WX433,WX1004);
  not NOT_142(WX437,WX1004);
  not NOT_143(WX439,WX430);
  not NOT_144(WX440,WX439);
  not NOT_145(WX443,WX1003);
  not NOT_146(WX447,WX1004);
  not NOT_147(WX451,WX1004);
  not NOT_148(WX453,WX444);
  not NOT_149(WX454,WX453);
  not NOT_150(WX457,WX1003);
  not NOT_151(WX461,WX1004);
  not NOT_152(WX465,WX1004);
  not NOT_153(WX467,WX458);
  not NOT_154(WX468,WX467);
  not NOT_155(WX471,WX1003);
  not NOT_156(WX475,WX1004);
  not NOT_157(WX479,WX1004);
  not NOT_158(WX481,WX472);
  not NOT_159(WX482,WX481);
  not NOT_160(WX483,WX485);
  not NOT_161(WX548,WX965);
  not NOT_162(WX549,WX967);
  not NOT_163(WX550,WX969);
  not NOT_164(WX551,WX971);
  not NOT_165(WX552,WX973);
  not NOT_166(WX553,WX975);
  not NOT_167(WX554,WX977);
  not NOT_168(WX555,WX979);
  not NOT_169(WX556,WX981);
  not NOT_170(WX557,WX983);
  not NOT_171(WX558,WX985);
  not NOT_172(WX559,WX987);
  not NOT_173(WX560,WX989);
  not NOT_174(WX561,WX991);
  not NOT_175(WX562,WX993);
  not NOT_176(WX563,WX995);
  not NOT_177(WX564,WX933);
  not NOT_178(WX565,WX935);
  not NOT_179(WX566,WX937);
  not NOT_180(WX567,WX939);
  not NOT_181(WX568,WX941);
  not NOT_182(WX569,WX943);
  not NOT_183(WX570,WX945);
  not NOT_184(WX571,WX947);
  not NOT_185(WX572,WX949);
  not NOT_186(WX573,WX951);
  not NOT_187(WX574,WX953);
  not NOT_188(WX575,WX955);
  not NOT_189(WX576,WX957);
  not NOT_190(WX577,WX959);
  not NOT_191(WX578,WX961);
  not NOT_192(WX579,WX963);
  not NOT_193(WX580,WX548);
  not NOT_194(WX581,WX549);
  not NOT_195(WX582,WX550);
  not NOT_196(WX583,WX551);
  not NOT_197(WX584,WX552);
  not NOT_198(WX585,WX553);
  not NOT_199(WX586,WX554);
  not NOT_200(WX587,WX555);
  not NOT_201(WX588,WX556);
  not NOT_202(WX589,WX557);
  not NOT_203(WX590,WX558);
  not NOT_204(WX591,WX559);
  not NOT_205(WX592,WX560);
  not NOT_206(WX593,WX561);
  not NOT_207(WX594,WX562);
  not NOT_208(WX595,WX563);
  not NOT_209(WX596,WX564);
  not NOT_210(WX597,WX565);
  not NOT_211(WX598,WX566);
  not NOT_212(WX599,WX567);
  not NOT_213(WX600,WX568);
  not NOT_214(WX601,WX569);
  not NOT_215(WX602,WX570);
  not NOT_216(WX603,WX571);
  not NOT_217(WX604,WX572);
  not NOT_218(WX605,WX573);
  not NOT_219(WX606,WX574);
  not NOT_220(WX607,WX575);
  not NOT_221(WX608,WX576);
  not NOT_222(WX609,WX577);
  not NOT_223(WX610,WX578);
  not NOT_224(WX611,WX579);
  not NOT_225(WX612,WX837);
  not NOT_226(WX613,WX839);
  not NOT_227(WX614,WX841);
  not NOT_228(WX615,WX843);
  not NOT_229(WX616,WX845);
  not NOT_230(WX617,WX847);
  not NOT_231(WX618,WX849);
  not NOT_232(WX619,WX851);
  not NOT_233(WX620,WX853);
  not NOT_234(WX621,WX855);
  not NOT_235(WX622,WX857);
  not NOT_236(WX623,WX859);
  not NOT_237(WX624,WX861);
  not NOT_238(WX625,WX863);
  not NOT_239(WX626,WX865);
  not NOT_240(WX627,WX867);
  not NOT_241(WX628,WX869);
  not NOT_242(WX629,WX871);
  not NOT_243(WX630,WX873);
  not NOT_244(WX631,WX875);
  not NOT_245(WX632,WX877);
  not NOT_246(WX633,WX879);
  not NOT_247(WX634,WX881);
  not NOT_248(WX635,WX883);
  not NOT_249(WX636,WX885);
  not NOT_250(WX637,WX887);
  not NOT_251(WX638,WX889);
  not NOT_252(WX639,WX891);
  not NOT_253(WX640,WX893);
  not NOT_254(WX641,WX895);
  not NOT_255(WX642,WX897);
  not NOT_256(WX643,WX899);
  not NOT_257(WX932,WX916);
  not NOT_258(WX933,WX932);
  not NOT_259(WX934,WX917);
  not NOT_260(WX935,WX934);
  not NOT_261(WX936,WX918);
  not NOT_262(WX937,WX936);
  not NOT_263(WX938,WX919);
  not NOT_264(WX939,WX938);
  not NOT_265(WX940,WX920);
  not NOT_266(WX941,WX940);
  not NOT_267(WX942,WX921);
  not NOT_268(WX943,WX942);
  not NOT_269(WX944,WX922);
  not NOT_270(WX945,WX944);
  not NOT_271(WX946,WX923);
  not NOT_272(WX947,WX946);
  not NOT_273(WX948,WX924);
  not NOT_274(WX949,WX948);
  not NOT_275(WX950,WX925);
  not NOT_276(WX951,WX950);
  not NOT_277(WX952,WX926);
  not NOT_278(WX953,WX952);
  not NOT_279(WX954,WX927);
  not NOT_280(WX955,WX954);
  not NOT_281(WX956,WX928);
  not NOT_282(WX957,WX956);
  not NOT_283(WX958,WX929);
  not NOT_284(WX959,WX958);
  not NOT_285(WX960,WX930);
  not NOT_286(WX961,WX960);
  not NOT_287(WX962,WX931);
  not NOT_288(WX963,WX962);
  not NOT_289(WX964,WX900);
  not NOT_290(WX965,WX964);
  not NOT_291(WX966,WX901);
  not NOT_292(WX967,WX966);
  not NOT_293(WX968,WX902);
  not NOT_294(WX969,WX968);
  not NOT_295(WX970,WX903);
  not NOT_296(WX971,WX970);
  not NOT_297(WX972,WX904);
  not NOT_298(WX973,WX972);
  not NOT_299(WX974,WX905);
  not NOT_300(WX975,WX974);
  not NOT_301(WX976,WX906);
  not NOT_302(WX977,WX976);
  not NOT_303(WX978,WX907);
  not NOT_304(WX979,WX978);
  not NOT_305(WX980,WX908);
  not NOT_306(WX981,WX980);
  not NOT_307(WX982,WX909);
  not NOT_308(WX983,WX982);
  not NOT_309(WX984,WX910);
  not NOT_310(WX985,WX984);
  not NOT_311(WX986,WX911);
  not NOT_312(WX987,WX986);
  not NOT_313(WX988,WX912);
  not NOT_314(WX989,WX988);
  not NOT_315(WX990,WX913);
  not NOT_316(WX991,WX990);
  not NOT_317(WX992,WX914);
  not NOT_318(WX993,WX992);
  not NOT_319(WX994,WX915);
  not NOT_320(WX995,WX994);
  not NOT_321(WX996,TM0);
  not NOT_322(WX997,TM0);
  not NOT_323(WX998,TM0);
  not NOT_324(WX999,TM1);
  not NOT_325(WX1000,TM1);
  not NOT_326(WX1001,WX1000);
  not NOT_327(WX1002,WX998);
  not NOT_328(WX1003,WX999);
  not NOT_329(WX1004,WX997);
  not NOT_330(WX1005,WX996);
  not NOT_331(WX1009,WX1005);
  not NOT_332(WX1011,WX1010);
  not NOT_333(DATA_9_31,WX1011);
  not NOT_334(WX1016,WX1005);
  not NOT_335(WX1018,WX1017);
  not NOT_336(DATA_9_30,WX1018);
  not NOT_337(WX1023,WX1005);
  not NOT_338(WX1025,WX1024);
  not NOT_339(DATA_9_29,WX1025);
  not NOT_340(WX1030,WX1005);
  not NOT_341(WX1032,WX1031);
  not NOT_342(DATA_9_28,WX1032);
  not NOT_343(WX1037,WX1005);
  not NOT_344(WX1039,WX1038);
  not NOT_345(DATA_9_27,WX1039);
  not NOT_346(WX1044,WX1005);
  not NOT_347(WX1046,WX1045);
  not NOT_348(DATA_9_26,WX1046);
  not NOT_349(WX1051,WX1005);
  not NOT_350(WX1053,WX1052);
  not NOT_351(DATA_9_25,WX1053);
  not NOT_352(WX1058,WX1005);
  not NOT_353(WX1060,WX1059);
  not NOT_354(DATA_9_24,WX1060);
  not NOT_355(WX1065,WX1005);
  not NOT_356(WX1067,WX1066);
  not NOT_357(DATA_9_23,WX1067);
  not NOT_358(WX1072,WX1005);
  not NOT_359(WX1074,WX1073);
  not NOT_360(DATA_9_22,WX1074);
  not NOT_361(WX1079,WX1005);
  not NOT_362(WX1081,WX1080);
  not NOT_363(DATA_9_21,WX1081);
  not NOT_364(WX1086,WX1005);
  not NOT_365(WX1088,WX1087);
  not NOT_366(DATA_9_20,WX1088);
  not NOT_367(WX1093,WX1005);
  not NOT_368(WX1095,WX1094);
  not NOT_369(DATA_9_19,WX1095);
  not NOT_370(WX1100,WX1005);
  not NOT_371(WX1102,WX1101);
  not NOT_372(DATA_9_18,WX1102);
  not NOT_373(WX1107,WX1005);
  not NOT_374(WX1109,WX1108);
  not NOT_375(DATA_9_17,WX1109);
  not NOT_376(WX1114,WX1005);
  not NOT_377(WX1116,WX1115);
  not NOT_378(DATA_9_16,WX1116);
  not NOT_379(WX1121,WX1005);
  not NOT_380(WX1123,WX1122);
  not NOT_381(DATA_9_15,WX1123);
  not NOT_382(WX1128,WX1005);
  not NOT_383(WX1130,WX1129);
  not NOT_384(DATA_9_14,WX1130);
  not NOT_385(WX1135,WX1005);
  not NOT_386(WX1137,WX1136);
  not NOT_387(DATA_9_13,WX1137);
  not NOT_388(WX1142,WX1005);
  not NOT_389(WX1144,WX1143);
  not NOT_390(DATA_9_12,WX1144);
  not NOT_391(WX1149,WX1005);
  not NOT_392(WX1151,WX1150);
  not NOT_393(DATA_9_11,WX1151);
  not NOT_394(WX1156,WX1005);
  not NOT_395(WX1158,WX1157);
  not NOT_396(DATA_9_10,WX1158);
  not NOT_397(WX1163,WX1005);
  not NOT_398(WX1165,WX1164);
  not NOT_399(DATA_9_9,WX1165);
  not NOT_400(WX1170,WX1005);
  not NOT_401(WX1172,WX1171);
  not NOT_402(DATA_9_8,WX1172);
  not NOT_403(WX1177,WX1005);
  not NOT_404(WX1179,WX1178);
  not NOT_405(DATA_9_7,WX1179);
  not NOT_406(WX1184,WX1005);
  not NOT_407(WX1186,WX1185);
  not NOT_408(DATA_9_6,WX1186);
  not NOT_409(WX1191,WX1005);
  not NOT_410(WX1193,WX1192);
  not NOT_411(DATA_9_5,WX1193);
  not NOT_412(WX1198,WX1005);
  not NOT_413(WX1200,WX1199);
  not NOT_414(DATA_9_4,WX1200);
  not NOT_415(WX1205,WX1005);
  not NOT_416(WX1207,WX1206);
  not NOT_417(DATA_9_3,WX1207);
  not NOT_418(WX1212,WX1005);
  not NOT_419(WX1214,WX1213);
  not NOT_420(DATA_9_2,WX1214);
  not NOT_421(WX1219,WX1005);
  not NOT_422(WX1221,WX1220);
  not NOT_423(DATA_9_1,WX1221);
  not NOT_424(WX1226,WX1005);
  not NOT_425(WX1228,WX1227);
  not NOT_426(DATA_9_0,WX1228);
  not NOT_427(WX1230,RESET);
  not NOT_428(WX1263,WX1230);
  not NOT_429(WX1330,WX2296);
  not NOT_430(WX1334,WX2297);
  not NOT_431(WX1338,WX2297);
  not NOT_432(WX1340,WX1331);
  not NOT_433(WX1341,WX1340);
  not NOT_434(WX1344,WX2296);
  not NOT_435(WX1348,WX2297);
  not NOT_436(WX1352,WX2297);
  not NOT_437(WX1354,WX1345);
  not NOT_438(WX1355,WX1354);
  not NOT_439(WX1358,WX2296);
  not NOT_440(WX1362,WX2297);
  not NOT_441(WX1366,WX2297);
  not NOT_442(WX1368,WX1359);
  not NOT_443(WX1369,WX1368);
  not NOT_444(WX1372,WX2296);
  not NOT_445(WX1376,WX2297);
  not NOT_446(WX1380,WX2297);
  not NOT_447(WX1382,WX1373);
  not NOT_448(WX1383,WX1382);
  not NOT_449(WX1386,WX2296);
  not NOT_450(WX1390,WX2297);
  not NOT_451(WX1394,WX2297);
  not NOT_452(WX1396,WX1387);
  not NOT_453(WX1397,WX1396);
  not NOT_454(WX1400,WX2296);
  not NOT_455(WX1404,WX2297);
  not NOT_456(WX1408,WX2297);
  not NOT_457(WX1410,WX1401);
  not NOT_458(WX1411,WX1410);
  not NOT_459(WX1414,WX2296);
  not NOT_460(WX1418,WX2297);
  not NOT_461(WX1422,WX2297);
  not NOT_462(WX1424,WX1415);
  not NOT_463(WX1425,WX1424);
  not NOT_464(WX1428,WX2296);
  not NOT_465(WX1432,WX2297);
  not NOT_466(WX1436,WX2297);
  not NOT_467(WX1438,WX1429);
  not NOT_468(WX1439,WX1438);
  not NOT_469(WX1442,WX2296);
  not NOT_470(WX1446,WX2297);
  not NOT_471(WX1450,WX2297);
  not NOT_472(WX1452,WX1443);
  not NOT_473(WX1453,WX1452);
  not NOT_474(WX1456,WX2296);
  not NOT_475(WX1460,WX2297);
  not NOT_476(WX1464,WX2297);
  not NOT_477(WX1466,WX1457);
  not NOT_478(WX1467,WX1466);
  not NOT_479(WX1470,WX2296);
  not NOT_480(WX1474,WX2297);
  not NOT_481(WX1478,WX2297);
  not NOT_482(WX1480,WX1471);
  not NOT_483(WX1481,WX1480);
  not NOT_484(WX1484,WX2296);
  not NOT_485(WX1488,WX2297);
  not NOT_486(WX1492,WX2297);
  not NOT_487(WX1494,WX1485);
  not NOT_488(WX1495,WX1494);
  not NOT_489(WX1498,WX2296);
  not NOT_490(WX1502,WX2297);
  not NOT_491(WX1506,WX2297);
  not NOT_492(WX1508,WX1499);
  not NOT_493(WX1509,WX1508);
  not NOT_494(WX1512,WX2296);
  not NOT_495(WX1516,WX2297);
  not NOT_496(WX1520,WX2297);
  not NOT_497(WX1522,WX1513);
  not NOT_498(WX1523,WX1522);
  not NOT_499(WX1526,WX2296);
  not NOT_500(WX1530,WX2297);
  not NOT_501(WX1534,WX2297);
  not NOT_502(WX1536,WX1527);
  not NOT_503(WX1537,WX1536);
  not NOT_504(WX1540,WX2296);
  not NOT_505(WX1544,WX2297);
  not NOT_506(WX1548,WX2297);
  not NOT_507(WX1550,WX1541);
  not NOT_508(WX1551,WX1550);
  not NOT_509(WX1554,WX2296);
  not NOT_510(WX1558,WX2297);
  not NOT_511(WX1562,WX2297);
  not NOT_512(WX1564,WX1555);
  not NOT_513(WX1565,WX1564);
  not NOT_514(WX1568,WX2296);
  not NOT_515(WX1572,WX2297);
  not NOT_516(WX1576,WX2297);
  not NOT_517(WX1578,WX1569);
  not NOT_518(WX1579,WX1578);
  not NOT_519(WX1582,WX2296);
  not NOT_520(WX1586,WX2297);
  not NOT_521(WX1590,WX2297);
  not NOT_522(WX1592,WX1583);
  not NOT_523(WX1593,WX1592);
  not NOT_524(WX1596,WX2296);
  not NOT_525(WX1600,WX2297);
  not NOT_526(WX1604,WX2297);
  not NOT_527(WX1606,WX1597);
  not NOT_528(WX1607,WX1606);
  not NOT_529(WX1610,WX2296);
  not NOT_530(WX1614,WX2297);
  not NOT_531(WX1618,WX2297);
  not NOT_532(WX1620,WX1611);
  not NOT_533(WX1621,WX1620);
  not NOT_534(WX1624,WX2296);
  not NOT_535(WX1628,WX2297);
  not NOT_536(WX1632,WX2297);
  not NOT_537(WX1634,WX1625);
  not NOT_538(WX1635,WX1634);
  not NOT_539(WX1638,WX2296);
  not NOT_540(WX1642,WX2297);
  not NOT_541(WX1646,WX2297);
  not NOT_542(WX1648,WX1639);
  not NOT_543(WX1649,WX1648);
  not NOT_544(WX1652,WX2296);
  not NOT_545(WX1656,WX2297);
  not NOT_546(WX1660,WX2297);
  not NOT_547(WX1662,WX1653);
  not NOT_548(WX1663,WX1662);
  not NOT_549(WX1666,WX2296);
  not NOT_550(WX1670,WX2297);
  not NOT_551(WX1674,WX2297);
  not NOT_552(WX1676,WX1667);
  not NOT_553(WX1677,WX1676);
  not NOT_554(WX1680,WX2296);
  not NOT_555(WX1684,WX2297);
  not NOT_556(WX1688,WX2297);
  not NOT_557(WX1690,WX1681);
  not NOT_558(WX1691,WX1690);
  not NOT_559(WX1694,WX2296);
  not NOT_560(WX1698,WX2297);
  not NOT_561(WX1702,WX2297);
  not NOT_562(WX1704,WX1695);
  not NOT_563(WX1705,WX1704);
  not NOT_564(WX1708,WX2296);
  not NOT_565(WX1712,WX2297);
  not NOT_566(WX1716,WX2297);
  not NOT_567(WX1718,WX1709);
  not NOT_568(WX1719,WX1718);
  not NOT_569(WX1722,WX2296);
  not NOT_570(WX1726,WX2297);
  not NOT_571(WX1730,WX2297);
  not NOT_572(WX1732,WX1723);
  not NOT_573(WX1733,WX1732);
  not NOT_574(WX1736,WX2296);
  not NOT_575(WX1740,WX2297);
  not NOT_576(WX1744,WX2297);
  not NOT_577(WX1746,WX1737);
  not NOT_578(WX1747,WX1746);
  not NOT_579(WX1750,WX2296);
  not NOT_580(WX1754,WX2297);
  not NOT_581(WX1758,WX2297);
  not NOT_582(WX1760,WX1751);
  not NOT_583(WX1761,WX1760);
  not NOT_584(WX1764,WX2296);
  not NOT_585(WX1768,WX2297);
  not NOT_586(WX1772,WX2297);
  not NOT_587(WX1774,WX1765);
  not NOT_588(WX1775,WX1774);
  not NOT_589(WX1776,WX1778);
  not NOT_590(WX1841,WX2258);
  not NOT_591(WX1842,WX2260);
  not NOT_592(WX1843,WX2262);
  not NOT_593(WX1844,WX2264);
  not NOT_594(WX1845,WX2266);
  not NOT_595(WX1846,WX2268);
  not NOT_596(WX1847,WX2270);
  not NOT_597(WX1848,WX2272);
  not NOT_598(WX1849,WX2274);
  not NOT_599(WX1850,WX2276);
  not NOT_600(WX1851,WX2278);
  not NOT_601(WX1852,WX2280);
  not NOT_602(WX1853,WX2282);
  not NOT_603(WX1854,WX2284);
  not NOT_604(WX1855,WX2286);
  not NOT_605(WX1856,WX2288);
  not NOT_606(WX1857,WX2226);
  not NOT_607(WX1858,WX2228);
  not NOT_608(WX1859,WX2230);
  not NOT_609(WX1860,WX2232);
  not NOT_610(WX1861,WX2234);
  not NOT_611(WX1862,WX2236);
  not NOT_612(WX1863,WX2238);
  not NOT_613(WX1864,WX2240);
  not NOT_614(WX1865,WX2242);
  not NOT_615(WX1866,WX2244);
  not NOT_616(WX1867,WX2246);
  not NOT_617(WX1868,WX2248);
  not NOT_618(WX1869,WX2250);
  not NOT_619(WX1870,WX2252);
  not NOT_620(WX1871,WX2254);
  not NOT_621(WX1872,WX2256);
  not NOT_622(WX1873,WX1841);
  not NOT_623(WX1874,WX1842);
  not NOT_624(WX1875,WX1843);
  not NOT_625(WX1876,WX1844);
  not NOT_626(WX1877,WX1845);
  not NOT_627(WX1878,WX1846);
  not NOT_628(WX1879,WX1847);
  not NOT_629(WX1880,WX1848);
  not NOT_630(WX1881,WX1849);
  not NOT_631(WX1882,WX1850);
  not NOT_632(WX1883,WX1851);
  not NOT_633(WX1884,WX1852);
  not NOT_634(WX1885,WX1853);
  not NOT_635(WX1886,WX1854);
  not NOT_636(WX1887,WX1855);
  not NOT_637(WX1888,WX1856);
  not NOT_638(WX1889,WX1857);
  not NOT_639(WX1890,WX1858);
  not NOT_640(WX1891,WX1859);
  not NOT_641(WX1892,WX1860);
  not NOT_642(WX1893,WX1861);
  not NOT_643(WX1894,WX1862);
  not NOT_644(WX1895,WX1863);
  not NOT_645(WX1896,WX1864);
  not NOT_646(WX1897,WX1865);
  not NOT_647(WX1898,WX1866);
  not NOT_648(WX1899,WX1867);
  not NOT_649(WX1900,WX1868);
  not NOT_650(WX1901,WX1869);
  not NOT_651(WX1902,WX1870);
  not NOT_652(WX1903,WX1871);
  not NOT_653(WX1904,WX1872);
  not NOT_654(WX1905,WX2130);
  not NOT_655(WX1906,WX2132);
  not NOT_656(WX1907,WX2134);
  not NOT_657(WX1908,WX2136);
  not NOT_658(WX1909,WX2138);
  not NOT_659(WX1910,WX2140);
  not NOT_660(WX1911,WX2142);
  not NOT_661(WX1912,WX2144);
  not NOT_662(WX1913,WX2146);
  not NOT_663(WX1914,WX2148);
  not NOT_664(WX1915,WX2150);
  not NOT_665(WX1916,WX2152);
  not NOT_666(WX1917,WX2154);
  not NOT_667(WX1918,WX2156);
  not NOT_668(WX1919,WX2158);
  not NOT_669(WX1920,WX2160);
  not NOT_670(WX1921,WX2162);
  not NOT_671(WX1922,WX2164);
  not NOT_672(WX1923,WX2166);
  not NOT_673(WX1924,WX2168);
  not NOT_674(WX1925,WX2170);
  not NOT_675(WX1926,WX2172);
  not NOT_676(WX1927,WX2174);
  not NOT_677(WX1928,WX2176);
  not NOT_678(WX1929,WX2178);
  not NOT_679(WX1930,WX2180);
  not NOT_680(WX1931,WX2182);
  not NOT_681(WX1932,WX2184);
  not NOT_682(WX1933,WX2186);
  not NOT_683(WX1934,WX2188);
  not NOT_684(WX1935,WX2190);
  not NOT_685(WX1936,WX2192);
  not NOT_686(WX2225,WX2209);
  not NOT_687(WX2226,WX2225);
  not NOT_688(WX2227,WX2210);
  not NOT_689(WX2228,WX2227);
  not NOT_690(WX2229,WX2211);
  not NOT_691(WX2230,WX2229);
  not NOT_692(WX2231,WX2212);
  not NOT_693(WX2232,WX2231);
  not NOT_694(WX2233,WX2213);
  not NOT_695(WX2234,WX2233);
  not NOT_696(WX2235,WX2214);
  not NOT_697(WX2236,WX2235);
  not NOT_698(WX2237,WX2215);
  not NOT_699(WX2238,WX2237);
  not NOT_700(WX2239,WX2216);
  not NOT_701(WX2240,WX2239);
  not NOT_702(WX2241,WX2217);
  not NOT_703(WX2242,WX2241);
  not NOT_704(WX2243,WX2218);
  not NOT_705(WX2244,WX2243);
  not NOT_706(WX2245,WX2219);
  not NOT_707(WX2246,WX2245);
  not NOT_708(WX2247,WX2220);
  not NOT_709(WX2248,WX2247);
  not NOT_710(WX2249,WX2221);
  not NOT_711(WX2250,WX2249);
  not NOT_712(WX2251,WX2222);
  not NOT_713(WX2252,WX2251);
  not NOT_714(WX2253,WX2223);
  not NOT_715(WX2254,WX2253);
  not NOT_716(WX2255,WX2224);
  not NOT_717(WX2256,WX2255);
  not NOT_718(WX2257,WX2193);
  not NOT_719(WX2258,WX2257);
  not NOT_720(WX2259,WX2194);
  not NOT_721(WX2260,WX2259);
  not NOT_722(WX2261,WX2195);
  not NOT_723(WX2262,WX2261);
  not NOT_724(WX2263,WX2196);
  not NOT_725(WX2264,WX2263);
  not NOT_726(WX2265,WX2197);
  not NOT_727(WX2266,WX2265);
  not NOT_728(WX2267,WX2198);
  not NOT_729(WX2268,WX2267);
  not NOT_730(WX2269,WX2199);
  not NOT_731(WX2270,WX2269);
  not NOT_732(WX2271,WX2200);
  not NOT_733(WX2272,WX2271);
  not NOT_734(WX2273,WX2201);
  not NOT_735(WX2274,WX2273);
  not NOT_736(WX2275,WX2202);
  not NOT_737(WX2276,WX2275);
  not NOT_738(WX2277,WX2203);
  not NOT_739(WX2278,WX2277);
  not NOT_740(WX2279,WX2204);
  not NOT_741(WX2280,WX2279);
  not NOT_742(WX2281,WX2205);
  not NOT_743(WX2282,WX2281);
  not NOT_744(WX2283,WX2206);
  not NOT_745(WX2284,WX2283);
  not NOT_746(WX2285,WX2207);
  not NOT_747(WX2286,WX2285);
  not NOT_748(WX2287,WX2208);
  not NOT_749(WX2288,WX2287);
  not NOT_750(WX2289,TM0);
  not NOT_751(WX2290,TM0);
  not NOT_752(WX2291,TM0);
  not NOT_753(WX2292,TM1);
  not NOT_754(WX2293,TM1);
  not NOT_755(WX2294,WX2293);
  not NOT_756(WX2295,WX2291);
  not NOT_757(WX2296,WX2292);
  not NOT_758(WX2297,WX2290);
  not NOT_759(WX2298,WX2289);
  not NOT_760(WX2302,WX2298);
  not NOT_761(WX2304,WX2303);
  not NOT_762(WX2305,WX2304);
  not NOT_763(WX2309,WX2298);
  not NOT_764(WX2311,WX2310);
  not NOT_765(WX2312,WX2311);
  not NOT_766(WX2316,WX2298);
  not NOT_767(WX2318,WX2317);
  not NOT_768(WX2319,WX2318);
  not NOT_769(WX2323,WX2298);
  not NOT_770(WX2325,WX2324);
  not NOT_771(WX2326,WX2325);
  not NOT_772(WX2330,WX2298);
  not NOT_773(WX2332,WX2331);
  not NOT_774(WX2333,WX2332);
  not NOT_775(WX2337,WX2298);
  not NOT_776(WX2339,WX2338);
  not NOT_777(WX2340,WX2339);
  not NOT_778(WX2344,WX2298);
  not NOT_779(WX2346,WX2345);
  not NOT_780(WX2347,WX2346);
  not NOT_781(WX2351,WX2298);
  not NOT_782(WX2353,WX2352);
  not NOT_783(WX2354,WX2353);
  not NOT_784(WX2358,WX2298);
  not NOT_785(WX2360,WX2359);
  not NOT_786(WX2361,WX2360);
  not NOT_787(WX2365,WX2298);
  not NOT_788(WX2367,WX2366);
  not NOT_789(WX2368,WX2367);
  not NOT_790(WX2372,WX2298);
  not NOT_791(WX2374,WX2373);
  not NOT_792(WX2375,WX2374);
  not NOT_793(WX2379,WX2298);
  not NOT_794(WX2381,WX2380);
  not NOT_795(WX2382,WX2381);
  not NOT_796(WX2386,WX2298);
  not NOT_797(WX2388,WX2387);
  not NOT_798(WX2389,WX2388);
  not NOT_799(WX2393,WX2298);
  not NOT_800(WX2395,WX2394);
  not NOT_801(WX2396,WX2395);
  not NOT_802(WX2400,WX2298);
  not NOT_803(WX2402,WX2401);
  not NOT_804(WX2403,WX2402);
  not NOT_805(WX2407,WX2298);
  not NOT_806(WX2409,WX2408);
  not NOT_807(WX2410,WX2409);
  not NOT_808(WX2414,WX2298);
  not NOT_809(WX2416,WX2415);
  not NOT_810(WX2417,WX2416);
  not NOT_811(WX2421,WX2298);
  not NOT_812(WX2423,WX2422);
  not NOT_813(WX2424,WX2423);
  not NOT_814(WX2428,WX2298);
  not NOT_815(WX2430,WX2429);
  not NOT_816(WX2431,WX2430);
  not NOT_817(WX2435,WX2298);
  not NOT_818(WX2437,WX2436);
  not NOT_819(WX2438,WX2437);
  not NOT_820(WX2442,WX2298);
  not NOT_821(WX2444,WX2443);
  not NOT_822(WX2445,WX2444);
  not NOT_823(WX2449,WX2298);
  not NOT_824(WX2451,WX2450);
  not NOT_825(WX2452,WX2451);
  not NOT_826(WX2456,WX2298);
  not NOT_827(WX2458,WX2457);
  not NOT_828(WX2459,WX2458);
  not NOT_829(WX2463,WX2298);
  not NOT_830(WX2465,WX2464);
  not NOT_831(WX2466,WX2465);
  not NOT_832(WX2470,WX2298);
  not NOT_833(WX2472,WX2471);
  not NOT_834(WX2473,WX2472);
  not NOT_835(WX2477,WX2298);
  not NOT_836(WX2479,WX2478);
  not NOT_837(WX2480,WX2479);
  not NOT_838(WX2484,WX2298);
  not NOT_839(WX2486,WX2485);
  not NOT_840(WX2487,WX2486);
  not NOT_841(WX2491,WX2298);
  not NOT_842(WX2493,WX2492);
  not NOT_843(WX2494,WX2493);
  not NOT_844(WX2498,WX2298);
  not NOT_845(WX2500,WX2499);
  not NOT_846(WX2501,WX2500);
  not NOT_847(WX2505,WX2298);
  not NOT_848(WX2507,WX2506);
  not NOT_849(WX2508,WX2507);
  not NOT_850(WX2512,WX2298);
  not NOT_851(WX2514,WX2513);
  not NOT_852(WX2515,WX2514);
  not NOT_853(WX2519,WX2298);
  not NOT_854(WX2521,WX2520);
  not NOT_855(WX2522,WX2521);
  not NOT_856(WX2523,RESET);
  not NOT_857(WX2556,WX2523);
  not NOT_858(WX2623,WX3589);
  not NOT_859(WX2627,WX3590);
  not NOT_860(WX2631,WX3590);
  not NOT_861(WX2633,WX2624);
  not NOT_862(WX2634,WX2633);
  not NOT_863(WX2637,WX3589);
  not NOT_864(WX2641,WX3590);
  not NOT_865(WX2645,WX3590);
  not NOT_866(WX2647,WX2638);
  not NOT_867(WX2648,WX2647);
  not NOT_868(WX2651,WX3589);
  not NOT_869(WX2655,WX3590);
  not NOT_870(WX2659,WX3590);
  not NOT_871(WX2661,WX2652);
  not NOT_872(WX2662,WX2661);
  not NOT_873(WX2665,WX3589);
  not NOT_874(WX2669,WX3590);
  not NOT_875(WX2673,WX3590);
  not NOT_876(WX2675,WX2666);
  not NOT_877(WX2676,WX2675);
  not NOT_878(WX2679,WX3589);
  not NOT_879(WX2683,WX3590);
  not NOT_880(WX2687,WX3590);
  not NOT_881(WX2689,WX2680);
  not NOT_882(WX2690,WX2689);
  not NOT_883(WX2693,WX3589);
  not NOT_884(WX2697,WX3590);
  not NOT_885(WX2701,WX3590);
  not NOT_886(WX2703,WX2694);
  not NOT_887(WX2704,WX2703);
  not NOT_888(WX2707,WX3589);
  not NOT_889(WX2711,WX3590);
  not NOT_890(WX2715,WX3590);
  not NOT_891(WX2717,WX2708);
  not NOT_892(WX2718,WX2717);
  not NOT_893(WX2721,WX3589);
  not NOT_894(WX2725,WX3590);
  not NOT_895(WX2729,WX3590);
  not NOT_896(WX2731,WX2722);
  not NOT_897(WX2732,WX2731);
  not NOT_898(WX2735,WX3589);
  not NOT_899(WX2739,WX3590);
  not NOT_900(WX2743,WX3590);
  not NOT_901(WX2745,WX2736);
  not NOT_902(WX2746,WX2745);
  not NOT_903(WX2749,WX3589);
  not NOT_904(WX2753,WX3590);
  not NOT_905(WX2757,WX3590);
  not NOT_906(WX2759,WX2750);
  not NOT_907(WX2760,WX2759);
  not NOT_908(WX2763,WX3589);
  not NOT_909(WX2767,WX3590);
  not NOT_910(WX2771,WX3590);
  not NOT_911(WX2773,WX2764);
  not NOT_912(WX2774,WX2773);
  not NOT_913(WX2777,WX3589);
  not NOT_914(WX2781,WX3590);
  not NOT_915(WX2785,WX3590);
  not NOT_916(WX2787,WX2778);
  not NOT_917(WX2788,WX2787);
  not NOT_918(WX2791,WX3589);
  not NOT_919(WX2795,WX3590);
  not NOT_920(WX2799,WX3590);
  not NOT_921(WX2801,WX2792);
  not NOT_922(WX2802,WX2801);
  not NOT_923(WX2805,WX3589);
  not NOT_924(WX2809,WX3590);
  not NOT_925(WX2813,WX3590);
  not NOT_926(WX2815,WX2806);
  not NOT_927(WX2816,WX2815);
  not NOT_928(WX2819,WX3589);
  not NOT_929(WX2823,WX3590);
  not NOT_930(WX2827,WX3590);
  not NOT_931(WX2829,WX2820);
  not NOT_932(WX2830,WX2829);
  not NOT_933(WX2833,WX3589);
  not NOT_934(WX2837,WX3590);
  not NOT_935(WX2841,WX3590);
  not NOT_936(WX2843,WX2834);
  not NOT_937(WX2844,WX2843);
  not NOT_938(WX2847,WX3589);
  not NOT_939(WX2851,WX3590);
  not NOT_940(WX2855,WX3590);
  not NOT_941(WX2857,WX2848);
  not NOT_942(WX2858,WX2857);
  not NOT_943(WX2861,WX3589);
  not NOT_944(WX2865,WX3590);
  not NOT_945(WX2869,WX3590);
  not NOT_946(WX2871,WX2862);
  not NOT_947(WX2872,WX2871);
  not NOT_948(WX2875,WX3589);
  not NOT_949(WX2879,WX3590);
  not NOT_950(WX2883,WX3590);
  not NOT_951(WX2885,WX2876);
  not NOT_952(WX2886,WX2885);
  not NOT_953(WX2889,WX3589);
  not NOT_954(WX2893,WX3590);
  not NOT_955(WX2897,WX3590);
  not NOT_956(WX2899,WX2890);
  not NOT_957(WX2900,WX2899);
  not NOT_958(WX2903,WX3589);
  not NOT_959(WX2907,WX3590);
  not NOT_960(WX2911,WX3590);
  not NOT_961(WX2913,WX2904);
  not NOT_962(WX2914,WX2913);
  not NOT_963(WX2917,WX3589);
  not NOT_964(WX2921,WX3590);
  not NOT_965(WX2925,WX3590);
  not NOT_966(WX2927,WX2918);
  not NOT_967(WX2928,WX2927);
  not NOT_968(WX2931,WX3589);
  not NOT_969(WX2935,WX3590);
  not NOT_970(WX2939,WX3590);
  not NOT_971(WX2941,WX2932);
  not NOT_972(WX2942,WX2941);
  not NOT_973(WX2945,WX3589);
  not NOT_974(WX2949,WX3590);
  not NOT_975(WX2953,WX3590);
  not NOT_976(WX2955,WX2946);
  not NOT_977(WX2956,WX2955);
  not NOT_978(WX2959,WX3589);
  not NOT_979(WX2963,WX3590);
  not NOT_980(WX2967,WX3590);
  not NOT_981(WX2969,WX2960);
  not NOT_982(WX2970,WX2969);
  not NOT_983(WX2973,WX3589);
  not NOT_984(WX2977,WX3590);
  not NOT_985(WX2981,WX3590);
  not NOT_986(WX2983,WX2974);
  not NOT_987(WX2984,WX2983);
  not NOT_988(WX2987,WX3589);
  not NOT_989(WX2991,WX3590);
  not NOT_990(WX2995,WX3590);
  not NOT_991(WX2997,WX2988);
  not NOT_992(WX2998,WX2997);
  not NOT_993(WX3001,WX3589);
  not NOT_994(WX3005,WX3590);
  not NOT_995(WX3009,WX3590);
  not NOT_996(WX3011,WX3002);
  not NOT_997(WX3012,WX3011);
  not NOT_998(WX3015,WX3589);
  not NOT_999(WX3019,WX3590);
  not NOT_1000(WX3023,WX3590);
  not NOT_1001(WX3025,WX3016);
  not NOT_1002(WX3026,WX3025);
  not NOT_1003(WX3029,WX3589);
  not NOT_1004(WX3033,WX3590);
  not NOT_1005(WX3037,WX3590);
  not NOT_1006(WX3039,WX3030);
  not NOT_1007(WX3040,WX3039);
  not NOT_1008(WX3043,WX3589);
  not NOT_1009(WX3047,WX3590);
  not NOT_1010(WX3051,WX3590);
  not NOT_1011(WX3053,WX3044);
  not NOT_1012(WX3054,WX3053);
  not NOT_1013(WX3057,WX3589);
  not NOT_1014(WX3061,WX3590);
  not NOT_1015(WX3065,WX3590);
  not NOT_1016(WX3067,WX3058);
  not NOT_1017(WX3068,WX3067);
  not NOT_1018(WX3069,WX3071);
  not NOT_1019(WX3134,WX3551);
  not NOT_1020(WX3135,WX3553);
  not NOT_1021(WX3136,WX3555);
  not NOT_1022(WX3137,WX3557);
  not NOT_1023(WX3138,WX3559);
  not NOT_1024(WX3139,WX3561);
  not NOT_1025(WX3140,WX3563);
  not NOT_1026(WX3141,WX3565);
  not NOT_1027(WX3142,WX3567);
  not NOT_1028(WX3143,WX3569);
  not NOT_1029(WX3144,WX3571);
  not NOT_1030(WX3145,WX3573);
  not NOT_1031(WX3146,WX3575);
  not NOT_1032(WX3147,WX3577);
  not NOT_1033(WX3148,WX3579);
  not NOT_1034(WX3149,WX3581);
  not NOT_1035(WX3150,WX3519);
  not NOT_1036(WX3151,WX3521);
  not NOT_1037(WX3152,WX3523);
  not NOT_1038(WX3153,WX3525);
  not NOT_1039(WX3154,WX3527);
  not NOT_1040(WX3155,WX3529);
  not NOT_1041(WX3156,WX3531);
  not NOT_1042(WX3157,WX3533);
  not NOT_1043(WX3158,WX3535);
  not NOT_1044(WX3159,WX3537);
  not NOT_1045(WX3160,WX3539);
  not NOT_1046(WX3161,WX3541);
  not NOT_1047(WX3162,WX3543);
  not NOT_1048(WX3163,WX3545);
  not NOT_1049(WX3164,WX3547);
  not NOT_1050(WX3165,WX3549);
  not NOT_1051(WX3166,WX3134);
  not NOT_1052(WX3167,WX3135);
  not NOT_1053(WX3168,WX3136);
  not NOT_1054(WX3169,WX3137);
  not NOT_1055(WX3170,WX3138);
  not NOT_1056(WX3171,WX3139);
  not NOT_1057(WX3172,WX3140);
  not NOT_1058(WX3173,WX3141);
  not NOT_1059(WX3174,WX3142);
  not NOT_1060(WX3175,WX3143);
  not NOT_1061(WX3176,WX3144);
  not NOT_1062(WX3177,WX3145);
  not NOT_1063(WX3178,WX3146);
  not NOT_1064(WX3179,WX3147);
  not NOT_1065(WX3180,WX3148);
  not NOT_1066(WX3181,WX3149);
  not NOT_1067(WX3182,WX3150);
  not NOT_1068(WX3183,WX3151);
  not NOT_1069(WX3184,WX3152);
  not NOT_1070(WX3185,WX3153);
  not NOT_1071(WX3186,WX3154);
  not NOT_1072(WX3187,WX3155);
  not NOT_1073(WX3188,WX3156);
  not NOT_1074(WX3189,WX3157);
  not NOT_1075(WX3190,WX3158);
  not NOT_1076(WX3191,WX3159);
  not NOT_1077(WX3192,WX3160);
  not NOT_1078(WX3193,WX3161);
  not NOT_1079(WX3194,WX3162);
  not NOT_1080(WX3195,WX3163);
  not NOT_1081(WX3196,WX3164);
  not NOT_1082(WX3197,WX3165);
  not NOT_1083(WX3198,WX3423);
  not NOT_1084(WX3199,WX3425);
  not NOT_1085(WX3200,WX3427);
  not NOT_1086(WX3201,WX3429);
  not NOT_1087(WX3202,WX3431);
  not NOT_1088(WX3203,WX3433);
  not NOT_1089(WX3204,WX3435);
  not NOT_1090(WX3205,WX3437);
  not NOT_1091(WX3206,WX3439);
  not NOT_1092(WX3207,WX3441);
  not NOT_1093(WX3208,WX3443);
  not NOT_1094(WX3209,WX3445);
  not NOT_1095(WX3210,WX3447);
  not NOT_1096(WX3211,WX3449);
  not NOT_1097(WX3212,WX3451);
  not NOT_1098(WX3213,WX3453);
  not NOT_1099(WX3214,WX3455);
  not NOT_1100(WX3215,WX3457);
  not NOT_1101(WX3216,WX3459);
  not NOT_1102(WX3217,WX3461);
  not NOT_1103(WX3218,WX3463);
  not NOT_1104(WX3219,WX3465);
  not NOT_1105(WX3220,WX3467);
  not NOT_1106(WX3221,WX3469);
  not NOT_1107(WX3222,WX3471);
  not NOT_1108(WX3223,WX3473);
  not NOT_1109(WX3224,WX3475);
  not NOT_1110(WX3225,WX3477);
  not NOT_1111(WX3226,WX3479);
  not NOT_1112(WX3227,WX3481);
  not NOT_1113(WX3228,WX3483);
  not NOT_1114(WX3229,WX3485);
  not NOT_1115(WX3518,WX3502);
  not NOT_1116(WX3519,WX3518);
  not NOT_1117(WX3520,WX3503);
  not NOT_1118(WX3521,WX3520);
  not NOT_1119(WX3522,WX3504);
  not NOT_1120(WX3523,WX3522);
  not NOT_1121(WX3524,WX3505);
  not NOT_1122(WX3525,WX3524);
  not NOT_1123(WX3526,WX3506);
  not NOT_1124(WX3527,WX3526);
  not NOT_1125(WX3528,WX3507);
  not NOT_1126(WX3529,WX3528);
  not NOT_1127(WX3530,WX3508);
  not NOT_1128(WX3531,WX3530);
  not NOT_1129(WX3532,WX3509);
  not NOT_1130(WX3533,WX3532);
  not NOT_1131(WX3534,WX3510);
  not NOT_1132(WX3535,WX3534);
  not NOT_1133(WX3536,WX3511);
  not NOT_1134(WX3537,WX3536);
  not NOT_1135(WX3538,WX3512);
  not NOT_1136(WX3539,WX3538);
  not NOT_1137(WX3540,WX3513);
  not NOT_1138(WX3541,WX3540);
  not NOT_1139(WX3542,WX3514);
  not NOT_1140(WX3543,WX3542);
  not NOT_1141(WX3544,WX3515);
  not NOT_1142(WX3545,WX3544);
  not NOT_1143(WX3546,WX3516);
  not NOT_1144(WX3547,WX3546);
  not NOT_1145(WX3548,WX3517);
  not NOT_1146(WX3549,WX3548);
  not NOT_1147(WX3550,WX3486);
  not NOT_1148(WX3551,WX3550);
  not NOT_1149(WX3552,WX3487);
  not NOT_1150(WX3553,WX3552);
  not NOT_1151(WX3554,WX3488);
  not NOT_1152(WX3555,WX3554);
  not NOT_1153(WX3556,WX3489);
  not NOT_1154(WX3557,WX3556);
  not NOT_1155(WX3558,WX3490);
  not NOT_1156(WX3559,WX3558);
  not NOT_1157(WX3560,WX3491);
  not NOT_1158(WX3561,WX3560);
  not NOT_1159(WX3562,WX3492);
  not NOT_1160(WX3563,WX3562);
  not NOT_1161(WX3564,WX3493);
  not NOT_1162(WX3565,WX3564);
  not NOT_1163(WX3566,WX3494);
  not NOT_1164(WX3567,WX3566);
  not NOT_1165(WX3568,WX3495);
  not NOT_1166(WX3569,WX3568);
  not NOT_1167(WX3570,WX3496);
  not NOT_1168(WX3571,WX3570);
  not NOT_1169(WX3572,WX3497);
  not NOT_1170(WX3573,WX3572);
  not NOT_1171(WX3574,WX3498);
  not NOT_1172(WX3575,WX3574);
  not NOT_1173(WX3576,WX3499);
  not NOT_1174(WX3577,WX3576);
  not NOT_1175(WX3578,WX3500);
  not NOT_1176(WX3579,WX3578);
  not NOT_1177(WX3580,WX3501);
  not NOT_1178(WX3581,WX3580);
  not NOT_1179(WX3582,TM0);
  not NOT_1180(WX3583,TM0);
  not NOT_1181(WX3584,TM0);
  not NOT_1182(WX3585,TM1);
  not NOT_1183(WX3586,TM1);
  not NOT_1184(WX3587,WX3586);
  not NOT_1185(WX3588,WX3584);
  not NOT_1186(WX3589,WX3585);
  not NOT_1187(WX3590,WX3583);
  not NOT_1188(WX3591,WX3582);
  not NOT_1189(WX3595,WX3591);
  not NOT_1190(WX3597,WX3596);
  not NOT_1191(WX3598,WX3597);
  not NOT_1192(WX3602,WX3591);
  not NOT_1193(WX3604,WX3603);
  not NOT_1194(WX3605,WX3604);
  not NOT_1195(WX3609,WX3591);
  not NOT_1196(WX3611,WX3610);
  not NOT_1197(WX3612,WX3611);
  not NOT_1198(WX3616,WX3591);
  not NOT_1199(WX3618,WX3617);
  not NOT_1200(WX3619,WX3618);
  not NOT_1201(WX3623,WX3591);
  not NOT_1202(WX3625,WX3624);
  not NOT_1203(WX3626,WX3625);
  not NOT_1204(WX3630,WX3591);
  not NOT_1205(WX3632,WX3631);
  not NOT_1206(WX3633,WX3632);
  not NOT_1207(WX3637,WX3591);
  not NOT_1208(WX3639,WX3638);
  not NOT_1209(WX3640,WX3639);
  not NOT_1210(WX3644,WX3591);
  not NOT_1211(WX3646,WX3645);
  not NOT_1212(WX3647,WX3646);
  not NOT_1213(WX3651,WX3591);
  not NOT_1214(WX3653,WX3652);
  not NOT_1215(WX3654,WX3653);
  not NOT_1216(WX3658,WX3591);
  not NOT_1217(WX3660,WX3659);
  not NOT_1218(WX3661,WX3660);
  not NOT_1219(WX3665,WX3591);
  not NOT_1220(WX3667,WX3666);
  not NOT_1221(WX3668,WX3667);
  not NOT_1222(WX3672,WX3591);
  not NOT_1223(WX3674,WX3673);
  not NOT_1224(WX3675,WX3674);
  not NOT_1225(WX3679,WX3591);
  not NOT_1226(WX3681,WX3680);
  not NOT_1227(WX3682,WX3681);
  not NOT_1228(WX3686,WX3591);
  not NOT_1229(WX3688,WX3687);
  not NOT_1230(WX3689,WX3688);
  not NOT_1231(WX3693,WX3591);
  not NOT_1232(WX3695,WX3694);
  not NOT_1233(WX3696,WX3695);
  not NOT_1234(WX3700,WX3591);
  not NOT_1235(WX3702,WX3701);
  not NOT_1236(WX3703,WX3702);
  not NOT_1237(WX3707,WX3591);
  not NOT_1238(WX3709,WX3708);
  not NOT_1239(WX3710,WX3709);
  not NOT_1240(WX3714,WX3591);
  not NOT_1241(WX3716,WX3715);
  not NOT_1242(WX3717,WX3716);
  not NOT_1243(WX3721,WX3591);
  not NOT_1244(WX3723,WX3722);
  not NOT_1245(WX3724,WX3723);
  not NOT_1246(WX3728,WX3591);
  not NOT_1247(WX3730,WX3729);
  not NOT_1248(WX3731,WX3730);
  not NOT_1249(WX3735,WX3591);
  not NOT_1250(WX3737,WX3736);
  not NOT_1251(WX3738,WX3737);
  not NOT_1252(WX3742,WX3591);
  not NOT_1253(WX3744,WX3743);
  not NOT_1254(WX3745,WX3744);
  not NOT_1255(WX3749,WX3591);
  not NOT_1256(WX3751,WX3750);
  not NOT_1257(WX3752,WX3751);
  not NOT_1258(WX3756,WX3591);
  not NOT_1259(WX3758,WX3757);
  not NOT_1260(WX3759,WX3758);
  not NOT_1261(WX3763,WX3591);
  not NOT_1262(WX3765,WX3764);
  not NOT_1263(WX3766,WX3765);
  not NOT_1264(WX3770,WX3591);
  not NOT_1265(WX3772,WX3771);
  not NOT_1266(WX3773,WX3772);
  not NOT_1267(WX3777,WX3591);
  not NOT_1268(WX3779,WX3778);
  not NOT_1269(WX3780,WX3779);
  not NOT_1270(WX3784,WX3591);
  not NOT_1271(WX3786,WX3785);
  not NOT_1272(WX3787,WX3786);
  not NOT_1273(WX3791,WX3591);
  not NOT_1274(WX3793,WX3792);
  not NOT_1275(WX3794,WX3793);
  not NOT_1276(WX3798,WX3591);
  not NOT_1277(WX3800,WX3799);
  not NOT_1278(WX3801,WX3800);
  not NOT_1279(WX3805,WX3591);
  not NOT_1280(WX3807,WX3806);
  not NOT_1281(WX3808,WX3807);
  not NOT_1282(WX3812,WX3591);
  not NOT_1283(WX3814,WX3813);
  not NOT_1284(WX3815,WX3814);
  not NOT_1285(WX3816,RESET);
  not NOT_1286(WX3849,WX3816);
  not NOT_1287(WX3916,WX4882);
  not NOT_1288(WX3920,WX4883);
  not NOT_1289(WX3924,WX4883);
  not NOT_1290(WX3926,WX3917);
  not NOT_1291(WX3927,WX3926);
  not NOT_1292(WX3930,WX4882);
  not NOT_1293(WX3934,WX4883);
  not NOT_1294(WX3938,WX4883);
  not NOT_1295(WX3940,WX3931);
  not NOT_1296(WX3941,WX3940);
  not NOT_1297(WX3944,WX4882);
  not NOT_1298(WX3948,WX4883);
  not NOT_1299(WX3952,WX4883);
  not NOT_1300(WX3954,WX3945);
  not NOT_1301(WX3955,WX3954);
  not NOT_1302(WX3958,WX4882);
  not NOT_1303(WX3962,WX4883);
  not NOT_1304(WX3966,WX4883);
  not NOT_1305(WX3968,WX3959);
  not NOT_1306(WX3969,WX3968);
  not NOT_1307(WX3972,WX4882);
  not NOT_1308(WX3976,WX4883);
  not NOT_1309(WX3980,WX4883);
  not NOT_1310(WX3982,WX3973);
  not NOT_1311(WX3983,WX3982);
  not NOT_1312(WX3986,WX4882);
  not NOT_1313(WX3990,WX4883);
  not NOT_1314(WX3994,WX4883);
  not NOT_1315(WX3996,WX3987);
  not NOT_1316(WX3997,WX3996);
  not NOT_1317(WX4000,WX4882);
  not NOT_1318(WX4004,WX4883);
  not NOT_1319(WX4008,WX4883);
  not NOT_1320(WX4010,WX4001);
  not NOT_1321(WX4011,WX4010);
  not NOT_1322(WX4014,WX4882);
  not NOT_1323(WX4018,WX4883);
  not NOT_1324(WX4022,WX4883);
  not NOT_1325(WX4024,WX4015);
  not NOT_1326(WX4025,WX4024);
  not NOT_1327(WX4028,WX4882);
  not NOT_1328(WX4032,WX4883);
  not NOT_1329(WX4036,WX4883);
  not NOT_1330(WX4038,WX4029);
  not NOT_1331(WX4039,WX4038);
  not NOT_1332(WX4042,WX4882);
  not NOT_1333(WX4046,WX4883);
  not NOT_1334(WX4050,WX4883);
  not NOT_1335(WX4052,WX4043);
  not NOT_1336(WX4053,WX4052);
  not NOT_1337(WX4056,WX4882);
  not NOT_1338(WX4060,WX4883);
  not NOT_1339(WX4064,WX4883);
  not NOT_1340(WX4066,WX4057);
  not NOT_1341(WX4067,WX4066);
  not NOT_1342(WX4070,WX4882);
  not NOT_1343(WX4074,WX4883);
  not NOT_1344(WX4078,WX4883);
  not NOT_1345(WX4080,WX4071);
  not NOT_1346(WX4081,WX4080);
  not NOT_1347(WX4084,WX4882);
  not NOT_1348(WX4088,WX4883);
  not NOT_1349(WX4092,WX4883);
  not NOT_1350(WX4094,WX4085);
  not NOT_1351(WX4095,WX4094);
  not NOT_1352(WX4098,WX4882);
  not NOT_1353(WX4102,WX4883);
  not NOT_1354(WX4106,WX4883);
  not NOT_1355(WX4108,WX4099);
  not NOT_1356(WX4109,WX4108);
  not NOT_1357(WX4112,WX4882);
  not NOT_1358(WX4116,WX4883);
  not NOT_1359(WX4120,WX4883);
  not NOT_1360(WX4122,WX4113);
  not NOT_1361(WX4123,WX4122);
  not NOT_1362(WX4126,WX4882);
  not NOT_1363(WX4130,WX4883);
  not NOT_1364(WX4134,WX4883);
  not NOT_1365(WX4136,WX4127);
  not NOT_1366(WX4137,WX4136);
  not NOT_1367(WX4140,WX4882);
  not NOT_1368(WX4144,WX4883);
  not NOT_1369(WX4148,WX4883);
  not NOT_1370(WX4150,WX4141);
  not NOT_1371(WX4151,WX4150);
  not NOT_1372(WX4154,WX4882);
  not NOT_1373(WX4158,WX4883);
  not NOT_1374(WX4162,WX4883);
  not NOT_1375(WX4164,WX4155);
  not NOT_1376(WX4165,WX4164);
  not NOT_1377(WX4168,WX4882);
  not NOT_1378(WX4172,WX4883);
  not NOT_1379(WX4176,WX4883);
  not NOT_1380(WX4178,WX4169);
  not NOT_1381(WX4179,WX4178);
  not NOT_1382(WX4182,WX4882);
  not NOT_1383(WX4186,WX4883);
  not NOT_1384(WX4190,WX4883);
  not NOT_1385(WX4192,WX4183);
  not NOT_1386(WX4193,WX4192);
  not NOT_1387(WX4196,WX4882);
  not NOT_1388(WX4200,WX4883);
  not NOT_1389(WX4204,WX4883);
  not NOT_1390(WX4206,WX4197);
  not NOT_1391(WX4207,WX4206);
  not NOT_1392(WX4210,WX4882);
  not NOT_1393(WX4214,WX4883);
  not NOT_1394(WX4218,WX4883);
  not NOT_1395(WX4220,WX4211);
  not NOT_1396(WX4221,WX4220);
  not NOT_1397(WX4224,WX4882);
  not NOT_1398(WX4228,WX4883);
  not NOT_1399(WX4232,WX4883);
  not NOT_1400(WX4234,WX4225);
  not NOT_1401(WX4235,WX4234);
  not NOT_1402(WX4238,WX4882);
  not NOT_1403(WX4242,WX4883);
  not NOT_1404(WX4246,WX4883);
  not NOT_1405(WX4248,WX4239);
  not NOT_1406(WX4249,WX4248);
  not NOT_1407(WX4252,WX4882);
  not NOT_1408(WX4256,WX4883);
  not NOT_1409(WX4260,WX4883);
  not NOT_1410(WX4262,WX4253);
  not NOT_1411(WX4263,WX4262);
  not NOT_1412(WX4266,WX4882);
  not NOT_1413(WX4270,WX4883);
  not NOT_1414(WX4274,WX4883);
  not NOT_1415(WX4276,WX4267);
  not NOT_1416(WX4277,WX4276);
  not NOT_1417(WX4280,WX4882);
  not NOT_1418(WX4284,WX4883);
  not NOT_1419(WX4288,WX4883);
  not NOT_1420(WX4290,WX4281);
  not NOT_1421(WX4291,WX4290);
  not NOT_1422(WX4294,WX4882);
  not NOT_1423(WX4298,WX4883);
  not NOT_1424(WX4302,WX4883);
  not NOT_1425(WX4304,WX4295);
  not NOT_1426(WX4305,WX4304);
  not NOT_1427(WX4308,WX4882);
  not NOT_1428(WX4312,WX4883);
  not NOT_1429(WX4316,WX4883);
  not NOT_1430(WX4318,WX4309);
  not NOT_1431(WX4319,WX4318);
  not NOT_1432(WX4322,WX4882);
  not NOT_1433(WX4326,WX4883);
  not NOT_1434(WX4330,WX4883);
  not NOT_1435(WX4332,WX4323);
  not NOT_1436(WX4333,WX4332);
  not NOT_1437(WX4336,WX4882);
  not NOT_1438(WX4340,WX4883);
  not NOT_1439(WX4344,WX4883);
  not NOT_1440(WX4346,WX4337);
  not NOT_1441(WX4347,WX4346);
  not NOT_1442(WX4350,WX4882);
  not NOT_1443(WX4354,WX4883);
  not NOT_1444(WX4358,WX4883);
  not NOT_1445(WX4360,WX4351);
  not NOT_1446(WX4361,WX4360);
  not NOT_1447(WX4362,WX4364);
  not NOT_1448(WX4427,WX4844);
  not NOT_1449(WX4428,WX4846);
  not NOT_1450(WX4429,WX4848);
  not NOT_1451(WX4430,WX4850);
  not NOT_1452(WX4431,WX4852);
  not NOT_1453(WX4432,WX4854);
  not NOT_1454(WX4433,WX4856);
  not NOT_1455(WX4434,WX4858);
  not NOT_1456(WX4435,WX4860);
  not NOT_1457(WX4436,WX4862);
  not NOT_1458(WX4437,WX4864);
  not NOT_1459(WX4438,WX4866);
  not NOT_1460(WX4439,WX4868);
  not NOT_1461(WX4440,WX4870);
  not NOT_1462(WX4441,WX4872);
  not NOT_1463(WX4442,WX4874);
  not NOT_1464(WX4443,WX4812);
  not NOT_1465(WX4444,WX4814);
  not NOT_1466(WX4445,WX4816);
  not NOT_1467(WX4446,WX4818);
  not NOT_1468(WX4447,WX4820);
  not NOT_1469(WX4448,WX4822);
  not NOT_1470(WX4449,WX4824);
  not NOT_1471(WX4450,WX4826);
  not NOT_1472(WX4451,WX4828);
  not NOT_1473(WX4452,WX4830);
  not NOT_1474(WX4453,WX4832);
  not NOT_1475(WX4454,WX4834);
  not NOT_1476(WX4455,WX4836);
  not NOT_1477(WX4456,WX4838);
  not NOT_1478(WX4457,WX4840);
  not NOT_1479(WX4458,WX4842);
  not NOT_1480(WX4459,WX4427);
  not NOT_1481(WX4460,WX4428);
  not NOT_1482(WX4461,WX4429);
  not NOT_1483(WX4462,WX4430);
  not NOT_1484(WX4463,WX4431);
  not NOT_1485(WX4464,WX4432);
  not NOT_1486(WX4465,WX4433);
  not NOT_1487(WX4466,WX4434);
  not NOT_1488(WX4467,WX4435);
  not NOT_1489(WX4468,WX4436);
  not NOT_1490(WX4469,WX4437);
  not NOT_1491(WX4470,WX4438);
  not NOT_1492(WX4471,WX4439);
  not NOT_1493(WX4472,WX4440);
  not NOT_1494(WX4473,WX4441);
  not NOT_1495(WX4474,WX4442);
  not NOT_1496(WX4475,WX4443);
  not NOT_1497(WX4476,WX4444);
  not NOT_1498(WX4477,WX4445);
  not NOT_1499(WX4478,WX4446);
  not NOT_1500(WX4479,WX4447);
  not NOT_1501(WX4480,WX4448);
  not NOT_1502(WX4481,WX4449);
  not NOT_1503(WX4482,WX4450);
  not NOT_1504(WX4483,WX4451);
  not NOT_1505(WX4484,WX4452);
  not NOT_1506(WX4485,WX4453);
  not NOT_1507(WX4486,WX4454);
  not NOT_1508(WX4487,WX4455);
  not NOT_1509(WX4488,WX4456);
  not NOT_1510(WX4489,WX4457);
  not NOT_1511(WX4490,WX4458);
  not NOT_1512(WX4491,WX4716);
  not NOT_1513(WX4492,WX4718);
  not NOT_1514(WX4493,WX4720);
  not NOT_1515(WX4494,WX4722);
  not NOT_1516(WX4495,WX4724);
  not NOT_1517(WX4496,WX4726);
  not NOT_1518(WX4497,WX4728);
  not NOT_1519(WX4498,WX4730);
  not NOT_1520(WX4499,WX4732);
  not NOT_1521(WX4500,WX4734);
  not NOT_1522(WX4501,WX4736);
  not NOT_1523(WX4502,WX4738);
  not NOT_1524(WX4503,WX4740);
  not NOT_1525(WX4504,WX4742);
  not NOT_1526(WX4505,WX4744);
  not NOT_1527(WX4506,WX4746);
  not NOT_1528(WX4507,WX4748);
  not NOT_1529(WX4508,WX4750);
  not NOT_1530(WX4509,WX4752);
  not NOT_1531(WX4510,WX4754);
  not NOT_1532(WX4511,WX4756);
  not NOT_1533(WX4512,WX4758);
  not NOT_1534(WX4513,WX4760);
  not NOT_1535(WX4514,WX4762);
  not NOT_1536(WX4515,WX4764);
  not NOT_1537(WX4516,WX4766);
  not NOT_1538(WX4517,WX4768);
  not NOT_1539(WX4518,WX4770);
  not NOT_1540(WX4519,WX4772);
  not NOT_1541(WX4520,WX4774);
  not NOT_1542(WX4521,WX4776);
  not NOT_1543(WX4522,WX4778);
  not NOT_1544(WX4811,WX4795);
  not NOT_1545(WX4812,WX4811);
  not NOT_1546(WX4813,WX4796);
  not NOT_1547(WX4814,WX4813);
  not NOT_1548(WX4815,WX4797);
  not NOT_1549(WX4816,WX4815);
  not NOT_1550(WX4817,WX4798);
  not NOT_1551(WX4818,WX4817);
  not NOT_1552(WX4819,WX4799);
  not NOT_1553(WX4820,WX4819);
  not NOT_1554(WX4821,WX4800);
  not NOT_1555(WX4822,WX4821);
  not NOT_1556(WX4823,WX4801);
  not NOT_1557(WX4824,WX4823);
  not NOT_1558(WX4825,WX4802);
  not NOT_1559(WX4826,WX4825);
  not NOT_1560(WX4827,WX4803);
  not NOT_1561(WX4828,WX4827);
  not NOT_1562(WX4829,WX4804);
  not NOT_1563(WX4830,WX4829);
  not NOT_1564(WX4831,WX4805);
  not NOT_1565(WX4832,WX4831);
  not NOT_1566(WX4833,WX4806);
  not NOT_1567(WX4834,WX4833);
  not NOT_1568(WX4835,WX4807);
  not NOT_1569(WX4836,WX4835);
  not NOT_1570(WX4837,WX4808);
  not NOT_1571(WX4838,WX4837);
  not NOT_1572(WX4839,WX4809);
  not NOT_1573(WX4840,WX4839);
  not NOT_1574(WX4841,WX4810);
  not NOT_1575(WX4842,WX4841);
  not NOT_1576(WX4843,WX4779);
  not NOT_1577(WX4844,WX4843);
  not NOT_1578(WX4845,WX4780);
  not NOT_1579(WX4846,WX4845);
  not NOT_1580(WX4847,WX4781);
  not NOT_1581(WX4848,WX4847);
  not NOT_1582(WX4849,WX4782);
  not NOT_1583(WX4850,WX4849);
  not NOT_1584(WX4851,WX4783);
  not NOT_1585(WX4852,WX4851);
  not NOT_1586(WX4853,WX4784);
  not NOT_1587(WX4854,WX4853);
  not NOT_1588(WX4855,WX4785);
  not NOT_1589(WX4856,WX4855);
  not NOT_1590(WX4857,WX4786);
  not NOT_1591(WX4858,WX4857);
  not NOT_1592(WX4859,WX4787);
  not NOT_1593(WX4860,WX4859);
  not NOT_1594(WX4861,WX4788);
  not NOT_1595(WX4862,WX4861);
  not NOT_1596(WX4863,WX4789);
  not NOT_1597(WX4864,WX4863);
  not NOT_1598(WX4865,WX4790);
  not NOT_1599(WX4866,WX4865);
  not NOT_1600(WX4867,WX4791);
  not NOT_1601(WX4868,WX4867);
  not NOT_1602(WX4869,WX4792);
  not NOT_1603(WX4870,WX4869);
  not NOT_1604(WX4871,WX4793);
  not NOT_1605(WX4872,WX4871);
  not NOT_1606(WX4873,WX4794);
  not NOT_1607(WX4874,WX4873);
  not NOT_1608(WX4875,TM0);
  not NOT_1609(WX4876,TM0);
  not NOT_1610(WX4877,TM0);
  not NOT_1611(WX4878,TM1);
  not NOT_1612(WX4879,TM1);
  not NOT_1613(WX4880,WX4879);
  not NOT_1614(WX4881,WX4877);
  not NOT_1615(WX4882,WX4878);
  not NOT_1616(WX4883,WX4876);
  not NOT_1617(WX4884,WX4875);
  not NOT_1618(WX4888,WX4884);
  not NOT_1619(WX4890,WX4889);
  not NOT_1620(WX4891,WX4890);
  not NOT_1621(WX4895,WX4884);
  not NOT_1622(WX4897,WX4896);
  not NOT_1623(WX4898,WX4897);
  not NOT_1624(WX4902,WX4884);
  not NOT_1625(WX4904,WX4903);
  not NOT_1626(WX4905,WX4904);
  not NOT_1627(WX4909,WX4884);
  not NOT_1628(WX4911,WX4910);
  not NOT_1629(WX4912,WX4911);
  not NOT_1630(WX4916,WX4884);
  not NOT_1631(WX4918,WX4917);
  not NOT_1632(WX4919,WX4918);
  not NOT_1633(WX4923,WX4884);
  not NOT_1634(WX4925,WX4924);
  not NOT_1635(WX4926,WX4925);
  not NOT_1636(WX4930,WX4884);
  not NOT_1637(WX4932,WX4931);
  not NOT_1638(WX4933,WX4932);
  not NOT_1639(WX4937,WX4884);
  not NOT_1640(WX4939,WX4938);
  not NOT_1641(WX4940,WX4939);
  not NOT_1642(WX4944,WX4884);
  not NOT_1643(WX4946,WX4945);
  not NOT_1644(WX4947,WX4946);
  not NOT_1645(WX4951,WX4884);
  not NOT_1646(WX4953,WX4952);
  not NOT_1647(WX4954,WX4953);
  not NOT_1648(WX4958,WX4884);
  not NOT_1649(WX4960,WX4959);
  not NOT_1650(WX4961,WX4960);
  not NOT_1651(WX4965,WX4884);
  not NOT_1652(WX4967,WX4966);
  not NOT_1653(WX4968,WX4967);
  not NOT_1654(WX4972,WX4884);
  not NOT_1655(WX4974,WX4973);
  not NOT_1656(WX4975,WX4974);
  not NOT_1657(WX4979,WX4884);
  not NOT_1658(WX4981,WX4980);
  not NOT_1659(WX4982,WX4981);
  not NOT_1660(WX4986,WX4884);
  not NOT_1661(WX4988,WX4987);
  not NOT_1662(WX4989,WX4988);
  not NOT_1663(WX4993,WX4884);
  not NOT_1664(WX4995,WX4994);
  not NOT_1665(WX4996,WX4995);
  not NOT_1666(WX5000,WX4884);
  not NOT_1667(WX5002,WX5001);
  not NOT_1668(WX5003,WX5002);
  not NOT_1669(WX5007,WX4884);
  not NOT_1670(WX5009,WX5008);
  not NOT_1671(WX5010,WX5009);
  not NOT_1672(WX5014,WX4884);
  not NOT_1673(WX5016,WX5015);
  not NOT_1674(WX5017,WX5016);
  not NOT_1675(WX5021,WX4884);
  not NOT_1676(WX5023,WX5022);
  not NOT_1677(WX5024,WX5023);
  not NOT_1678(WX5028,WX4884);
  not NOT_1679(WX5030,WX5029);
  not NOT_1680(WX5031,WX5030);
  not NOT_1681(WX5035,WX4884);
  not NOT_1682(WX5037,WX5036);
  not NOT_1683(WX5038,WX5037);
  not NOT_1684(WX5042,WX4884);
  not NOT_1685(WX5044,WX5043);
  not NOT_1686(WX5045,WX5044);
  not NOT_1687(WX5049,WX4884);
  not NOT_1688(WX5051,WX5050);
  not NOT_1689(WX5052,WX5051);
  not NOT_1690(WX5056,WX4884);
  not NOT_1691(WX5058,WX5057);
  not NOT_1692(WX5059,WX5058);
  not NOT_1693(WX5063,WX4884);
  not NOT_1694(WX5065,WX5064);
  not NOT_1695(WX5066,WX5065);
  not NOT_1696(WX5070,WX4884);
  not NOT_1697(WX5072,WX5071);
  not NOT_1698(WX5073,WX5072);
  not NOT_1699(WX5077,WX4884);
  not NOT_1700(WX5079,WX5078);
  not NOT_1701(WX5080,WX5079);
  not NOT_1702(WX5084,WX4884);
  not NOT_1703(WX5086,WX5085);
  not NOT_1704(WX5087,WX5086);
  not NOT_1705(WX5091,WX4884);
  not NOT_1706(WX5093,WX5092);
  not NOT_1707(WX5094,WX5093);
  not NOT_1708(WX5098,WX4884);
  not NOT_1709(WX5100,WX5099);
  not NOT_1710(WX5101,WX5100);
  not NOT_1711(WX5105,WX4884);
  not NOT_1712(WX5107,WX5106);
  not NOT_1713(WX5108,WX5107);
  not NOT_1714(WX5109,RESET);
  not NOT_1715(WX5142,WX5109);
  not NOT_1716(WX5209,WX6175);
  not NOT_1717(WX5213,WX6176);
  not NOT_1718(WX5217,WX6176);
  not NOT_1719(WX5219,WX5210);
  not NOT_1720(WX5220,WX5219);
  not NOT_1721(WX5223,WX6175);
  not NOT_1722(WX5227,WX6176);
  not NOT_1723(WX5231,WX6176);
  not NOT_1724(WX5233,WX5224);
  not NOT_1725(WX5234,WX5233);
  not NOT_1726(WX5237,WX6175);
  not NOT_1727(WX5241,WX6176);
  not NOT_1728(WX5245,WX6176);
  not NOT_1729(WX5247,WX5238);
  not NOT_1730(WX5248,WX5247);
  not NOT_1731(WX5251,WX6175);
  not NOT_1732(WX5255,WX6176);
  not NOT_1733(WX5259,WX6176);
  not NOT_1734(WX5261,WX5252);
  not NOT_1735(WX5262,WX5261);
  not NOT_1736(WX5265,WX6175);
  not NOT_1737(WX5269,WX6176);
  not NOT_1738(WX5273,WX6176);
  not NOT_1739(WX5275,WX5266);
  not NOT_1740(WX5276,WX5275);
  not NOT_1741(WX5279,WX6175);
  not NOT_1742(WX5283,WX6176);
  not NOT_1743(WX5287,WX6176);
  not NOT_1744(WX5289,WX5280);
  not NOT_1745(WX5290,WX5289);
  not NOT_1746(WX5293,WX6175);
  not NOT_1747(WX5297,WX6176);
  not NOT_1748(WX5301,WX6176);
  not NOT_1749(WX5303,WX5294);
  not NOT_1750(WX5304,WX5303);
  not NOT_1751(WX5307,WX6175);
  not NOT_1752(WX5311,WX6176);
  not NOT_1753(WX5315,WX6176);
  not NOT_1754(WX5317,WX5308);
  not NOT_1755(WX5318,WX5317);
  not NOT_1756(WX5321,WX6175);
  not NOT_1757(WX5325,WX6176);
  not NOT_1758(WX5329,WX6176);
  not NOT_1759(WX5331,WX5322);
  not NOT_1760(WX5332,WX5331);
  not NOT_1761(WX5335,WX6175);
  not NOT_1762(WX5339,WX6176);
  not NOT_1763(WX5343,WX6176);
  not NOT_1764(WX5345,WX5336);
  not NOT_1765(WX5346,WX5345);
  not NOT_1766(WX5349,WX6175);
  not NOT_1767(WX5353,WX6176);
  not NOT_1768(WX5357,WX6176);
  not NOT_1769(WX5359,WX5350);
  not NOT_1770(WX5360,WX5359);
  not NOT_1771(WX5363,WX6175);
  not NOT_1772(WX5367,WX6176);
  not NOT_1773(WX5371,WX6176);
  not NOT_1774(WX5373,WX5364);
  not NOT_1775(WX5374,WX5373);
  not NOT_1776(WX5377,WX6175);
  not NOT_1777(WX5381,WX6176);
  not NOT_1778(WX5385,WX6176);
  not NOT_1779(WX5387,WX5378);
  not NOT_1780(WX5388,WX5387);
  not NOT_1781(WX5391,WX6175);
  not NOT_1782(WX5395,WX6176);
  not NOT_1783(WX5399,WX6176);
  not NOT_1784(WX5401,WX5392);
  not NOT_1785(WX5402,WX5401);
  not NOT_1786(WX5405,WX6175);
  not NOT_1787(WX5409,WX6176);
  not NOT_1788(WX5413,WX6176);
  not NOT_1789(WX5415,WX5406);
  not NOT_1790(WX5416,WX5415);
  not NOT_1791(WX5419,WX6175);
  not NOT_1792(WX5423,WX6176);
  not NOT_1793(WX5427,WX6176);
  not NOT_1794(WX5429,WX5420);
  not NOT_1795(WX5430,WX5429);
  not NOT_1796(WX5433,WX6175);
  not NOT_1797(WX5437,WX6176);
  not NOT_1798(WX5441,WX6176);
  not NOT_1799(WX5443,WX5434);
  not NOT_1800(WX5444,WX5443);
  not NOT_1801(WX5447,WX6175);
  not NOT_1802(WX5451,WX6176);
  not NOT_1803(WX5455,WX6176);
  not NOT_1804(WX5457,WX5448);
  not NOT_1805(WX5458,WX5457);
  not NOT_1806(WX5461,WX6175);
  not NOT_1807(WX5465,WX6176);
  not NOT_1808(WX5469,WX6176);
  not NOT_1809(WX5471,WX5462);
  not NOT_1810(WX5472,WX5471);
  not NOT_1811(WX5475,WX6175);
  not NOT_1812(WX5479,WX6176);
  not NOT_1813(WX5483,WX6176);
  not NOT_1814(WX5485,WX5476);
  not NOT_1815(WX5486,WX5485);
  not NOT_1816(WX5489,WX6175);
  not NOT_1817(WX5493,WX6176);
  not NOT_1818(WX5497,WX6176);
  not NOT_1819(WX5499,WX5490);
  not NOT_1820(WX5500,WX5499);
  not NOT_1821(WX5503,WX6175);
  not NOT_1822(WX5507,WX6176);
  not NOT_1823(WX5511,WX6176);
  not NOT_1824(WX5513,WX5504);
  not NOT_1825(WX5514,WX5513);
  not NOT_1826(WX5517,WX6175);
  not NOT_1827(WX5521,WX6176);
  not NOT_1828(WX5525,WX6176);
  not NOT_1829(WX5527,WX5518);
  not NOT_1830(WX5528,WX5527);
  not NOT_1831(WX5531,WX6175);
  not NOT_1832(WX5535,WX6176);
  not NOT_1833(WX5539,WX6176);
  not NOT_1834(WX5541,WX5532);
  not NOT_1835(WX5542,WX5541);
  not NOT_1836(WX5545,WX6175);
  not NOT_1837(WX5549,WX6176);
  not NOT_1838(WX5553,WX6176);
  not NOT_1839(WX5555,WX5546);
  not NOT_1840(WX5556,WX5555);
  not NOT_1841(WX5559,WX6175);
  not NOT_1842(WX5563,WX6176);
  not NOT_1843(WX5567,WX6176);
  not NOT_1844(WX5569,WX5560);
  not NOT_1845(WX5570,WX5569);
  not NOT_1846(WX5573,WX6175);
  not NOT_1847(WX5577,WX6176);
  not NOT_1848(WX5581,WX6176);
  not NOT_1849(WX5583,WX5574);
  not NOT_1850(WX5584,WX5583);
  not NOT_1851(WX5587,WX6175);
  not NOT_1852(WX5591,WX6176);
  not NOT_1853(WX5595,WX6176);
  not NOT_1854(WX5597,WX5588);
  not NOT_1855(WX5598,WX5597);
  not NOT_1856(WX5601,WX6175);
  not NOT_1857(WX5605,WX6176);
  not NOT_1858(WX5609,WX6176);
  not NOT_1859(WX5611,WX5602);
  not NOT_1860(WX5612,WX5611);
  not NOT_1861(WX5615,WX6175);
  not NOT_1862(WX5619,WX6176);
  not NOT_1863(WX5623,WX6176);
  not NOT_1864(WX5625,WX5616);
  not NOT_1865(WX5626,WX5625);
  not NOT_1866(WX5629,WX6175);
  not NOT_1867(WX5633,WX6176);
  not NOT_1868(WX5637,WX6176);
  not NOT_1869(WX5639,WX5630);
  not NOT_1870(WX5640,WX5639);
  not NOT_1871(WX5643,WX6175);
  not NOT_1872(WX5647,WX6176);
  not NOT_1873(WX5651,WX6176);
  not NOT_1874(WX5653,WX5644);
  not NOT_1875(WX5654,WX5653);
  not NOT_1876(WX5655,WX5657);
  not NOT_1877(WX5720,WX6137);
  not NOT_1878(WX5721,WX6139);
  not NOT_1879(WX5722,WX6141);
  not NOT_1880(WX5723,WX6143);
  not NOT_1881(WX5724,WX6145);
  not NOT_1882(WX5725,WX6147);
  not NOT_1883(WX5726,WX6149);
  not NOT_1884(WX5727,WX6151);
  not NOT_1885(WX5728,WX6153);
  not NOT_1886(WX5729,WX6155);
  not NOT_1887(WX5730,WX6157);
  not NOT_1888(WX5731,WX6159);
  not NOT_1889(WX5732,WX6161);
  not NOT_1890(WX5733,WX6163);
  not NOT_1891(WX5734,WX6165);
  not NOT_1892(WX5735,WX6167);
  not NOT_1893(WX5736,WX6105);
  not NOT_1894(WX5737,WX6107);
  not NOT_1895(WX5738,WX6109);
  not NOT_1896(WX5739,WX6111);
  not NOT_1897(WX5740,WX6113);
  not NOT_1898(WX5741,WX6115);
  not NOT_1899(WX5742,WX6117);
  not NOT_1900(WX5743,WX6119);
  not NOT_1901(WX5744,WX6121);
  not NOT_1902(WX5745,WX6123);
  not NOT_1903(WX5746,WX6125);
  not NOT_1904(WX5747,WX6127);
  not NOT_1905(WX5748,WX6129);
  not NOT_1906(WX5749,WX6131);
  not NOT_1907(WX5750,WX6133);
  not NOT_1908(WX5751,WX6135);
  not NOT_1909(WX5752,WX5720);
  not NOT_1910(WX5753,WX5721);
  not NOT_1911(WX5754,WX5722);
  not NOT_1912(WX5755,WX5723);
  not NOT_1913(WX5756,WX5724);
  not NOT_1914(WX5757,WX5725);
  not NOT_1915(WX5758,WX5726);
  not NOT_1916(WX5759,WX5727);
  not NOT_1917(WX5760,WX5728);
  not NOT_1918(WX5761,WX5729);
  not NOT_1919(WX5762,WX5730);
  not NOT_1920(WX5763,WX5731);
  not NOT_1921(WX5764,WX5732);
  not NOT_1922(WX5765,WX5733);
  not NOT_1923(WX5766,WX5734);
  not NOT_1924(WX5767,WX5735);
  not NOT_1925(WX5768,WX5736);
  not NOT_1926(WX5769,WX5737);
  not NOT_1927(WX5770,WX5738);
  not NOT_1928(WX5771,WX5739);
  not NOT_1929(WX5772,WX5740);
  not NOT_1930(WX5773,WX5741);
  not NOT_1931(WX5774,WX5742);
  not NOT_1932(WX5775,WX5743);
  not NOT_1933(WX5776,WX5744);
  not NOT_1934(WX5777,WX5745);
  not NOT_1935(WX5778,WX5746);
  not NOT_1936(WX5779,WX5747);
  not NOT_1937(WX5780,WX5748);
  not NOT_1938(WX5781,WX5749);
  not NOT_1939(WX5782,WX5750);
  not NOT_1940(WX5783,WX5751);
  not NOT_1941(WX5784,WX6009);
  not NOT_1942(WX5785,WX6011);
  not NOT_1943(WX5786,WX6013);
  not NOT_1944(WX5787,WX6015);
  not NOT_1945(WX5788,WX6017);
  not NOT_1946(WX5789,WX6019);
  not NOT_1947(WX5790,WX6021);
  not NOT_1948(WX5791,WX6023);
  not NOT_1949(WX5792,WX6025);
  not NOT_1950(WX5793,WX6027);
  not NOT_1951(WX5794,WX6029);
  not NOT_1952(WX5795,WX6031);
  not NOT_1953(WX5796,WX6033);
  not NOT_1954(WX5797,WX6035);
  not NOT_1955(WX5798,WX6037);
  not NOT_1956(WX5799,WX6039);
  not NOT_1957(WX5800,WX6041);
  not NOT_1958(WX5801,WX6043);
  not NOT_1959(WX5802,WX6045);
  not NOT_1960(WX5803,WX6047);
  not NOT_1961(WX5804,WX6049);
  not NOT_1962(WX5805,WX6051);
  not NOT_1963(WX5806,WX6053);
  not NOT_1964(WX5807,WX6055);
  not NOT_1965(WX5808,WX6057);
  not NOT_1966(WX5809,WX6059);
  not NOT_1967(WX5810,WX6061);
  not NOT_1968(WX5811,WX6063);
  not NOT_1969(WX5812,WX6065);
  not NOT_1970(WX5813,WX6067);
  not NOT_1971(WX5814,WX6069);
  not NOT_1972(WX5815,WX6071);
  not NOT_1973(WX6104,WX6088);
  not NOT_1974(WX6105,WX6104);
  not NOT_1975(WX6106,WX6089);
  not NOT_1976(WX6107,WX6106);
  not NOT_1977(WX6108,WX6090);
  not NOT_1978(WX6109,WX6108);
  not NOT_1979(WX6110,WX6091);
  not NOT_1980(WX6111,WX6110);
  not NOT_1981(WX6112,WX6092);
  not NOT_1982(WX6113,WX6112);
  not NOT_1983(WX6114,WX6093);
  not NOT_1984(WX6115,WX6114);
  not NOT_1985(WX6116,WX6094);
  not NOT_1986(WX6117,WX6116);
  not NOT_1987(WX6118,WX6095);
  not NOT_1988(WX6119,WX6118);
  not NOT_1989(WX6120,WX6096);
  not NOT_1990(WX6121,WX6120);
  not NOT_1991(WX6122,WX6097);
  not NOT_1992(WX6123,WX6122);
  not NOT_1993(WX6124,WX6098);
  not NOT_1994(WX6125,WX6124);
  not NOT_1995(WX6126,WX6099);
  not NOT_1996(WX6127,WX6126);
  not NOT_1997(WX6128,WX6100);
  not NOT_1998(WX6129,WX6128);
  not NOT_1999(WX6130,WX6101);
  not NOT_2000(WX6131,WX6130);
  not NOT_2001(WX6132,WX6102);
  not NOT_2002(WX6133,WX6132);
  not NOT_2003(WX6134,WX6103);
  not NOT_2004(WX6135,WX6134);
  not NOT_2005(WX6136,WX6072);
  not NOT_2006(WX6137,WX6136);
  not NOT_2007(WX6138,WX6073);
  not NOT_2008(WX6139,WX6138);
  not NOT_2009(WX6140,WX6074);
  not NOT_2010(WX6141,WX6140);
  not NOT_2011(WX6142,WX6075);
  not NOT_2012(WX6143,WX6142);
  not NOT_2013(WX6144,WX6076);
  not NOT_2014(WX6145,WX6144);
  not NOT_2015(WX6146,WX6077);
  not NOT_2016(WX6147,WX6146);
  not NOT_2017(WX6148,WX6078);
  not NOT_2018(WX6149,WX6148);
  not NOT_2019(WX6150,WX6079);
  not NOT_2020(WX6151,WX6150);
  not NOT_2021(WX6152,WX6080);
  not NOT_2022(WX6153,WX6152);
  not NOT_2023(WX6154,WX6081);
  not NOT_2024(WX6155,WX6154);
  not NOT_2025(WX6156,WX6082);
  not NOT_2026(WX6157,WX6156);
  not NOT_2027(WX6158,WX6083);
  not NOT_2028(WX6159,WX6158);
  not NOT_2029(WX6160,WX6084);
  not NOT_2030(WX6161,WX6160);
  not NOT_2031(WX6162,WX6085);
  not NOT_2032(WX6163,WX6162);
  not NOT_2033(WX6164,WX6086);
  not NOT_2034(WX6165,WX6164);
  not NOT_2035(WX6166,WX6087);
  not NOT_2036(WX6167,WX6166);
  not NOT_2037(WX6168,TM0);
  not NOT_2038(WX6169,TM0);
  not NOT_2039(WX6170,TM0);
  not NOT_2040(WX6171,TM1);
  not NOT_2041(WX6172,TM1);
  not NOT_2042(WX6173,WX6172);
  not NOT_2043(WX6174,WX6170);
  not NOT_2044(WX6175,WX6171);
  not NOT_2045(WX6176,WX6169);
  not NOT_2046(WX6177,WX6168);
  not NOT_2047(WX6181,WX6177);
  not NOT_2048(WX6183,WX6182);
  not NOT_2049(WX6184,WX6183);
  not NOT_2050(WX6188,WX6177);
  not NOT_2051(WX6190,WX6189);
  not NOT_2052(WX6191,WX6190);
  not NOT_2053(WX6195,WX6177);
  not NOT_2054(WX6197,WX6196);
  not NOT_2055(WX6198,WX6197);
  not NOT_2056(WX6202,WX6177);
  not NOT_2057(WX6204,WX6203);
  not NOT_2058(WX6205,WX6204);
  not NOT_2059(WX6209,WX6177);
  not NOT_2060(WX6211,WX6210);
  not NOT_2061(WX6212,WX6211);
  not NOT_2062(WX6216,WX6177);
  not NOT_2063(WX6218,WX6217);
  not NOT_2064(WX6219,WX6218);
  not NOT_2065(WX6223,WX6177);
  not NOT_2066(WX6225,WX6224);
  not NOT_2067(WX6226,WX6225);
  not NOT_2068(WX6230,WX6177);
  not NOT_2069(WX6232,WX6231);
  not NOT_2070(WX6233,WX6232);
  not NOT_2071(WX6237,WX6177);
  not NOT_2072(WX6239,WX6238);
  not NOT_2073(WX6240,WX6239);
  not NOT_2074(WX6244,WX6177);
  not NOT_2075(WX6246,WX6245);
  not NOT_2076(WX6247,WX6246);
  not NOT_2077(WX6251,WX6177);
  not NOT_2078(WX6253,WX6252);
  not NOT_2079(WX6254,WX6253);
  not NOT_2080(WX6258,WX6177);
  not NOT_2081(WX6260,WX6259);
  not NOT_2082(WX6261,WX6260);
  not NOT_2083(WX6265,WX6177);
  not NOT_2084(WX6267,WX6266);
  not NOT_2085(WX6268,WX6267);
  not NOT_2086(WX6272,WX6177);
  not NOT_2087(WX6274,WX6273);
  not NOT_2088(WX6275,WX6274);
  not NOT_2089(WX6279,WX6177);
  not NOT_2090(WX6281,WX6280);
  not NOT_2091(WX6282,WX6281);
  not NOT_2092(WX6286,WX6177);
  not NOT_2093(WX6288,WX6287);
  not NOT_2094(WX6289,WX6288);
  not NOT_2095(WX6293,WX6177);
  not NOT_2096(WX6295,WX6294);
  not NOT_2097(WX6296,WX6295);
  not NOT_2098(WX6300,WX6177);
  not NOT_2099(WX6302,WX6301);
  not NOT_2100(WX6303,WX6302);
  not NOT_2101(WX6307,WX6177);
  not NOT_2102(WX6309,WX6308);
  not NOT_2103(WX6310,WX6309);
  not NOT_2104(WX6314,WX6177);
  not NOT_2105(WX6316,WX6315);
  not NOT_2106(WX6317,WX6316);
  not NOT_2107(WX6321,WX6177);
  not NOT_2108(WX6323,WX6322);
  not NOT_2109(WX6324,WX6323);
  not NOT_2110(WX6328,WX6177);
  not NOT_2111(WX6330,WX6329);
  not NOT_2112(WX6331,WX6330);
  not NOT_2113(WX6335,WX6177);
  not NOT_2114(WX6337,WX6336);
  not NOT_2115(WX6338,WX6337);
  not NOT_2116(WX6342,WX6177);
  not NOT_2117(WX6344,WX6343);
  not NOT_2118(WX6345,WX6344);
  not NOT_2119(WX6349,WX6177);
  not NOT_2120(WX6351,WX6350);
  not NOT_2121(WX6352,WX6351);
  not NOT_2122(WX6356,WX6177);
  not NOT_2123(WX6358,WX6357);
  not NOT_2124(WX6359,WX6358);
  not NOT_2125(WX6363,WX6177);
  not NOT_2126(WX6365,WX6364);
  not NOT_2127(WX6366,WX6365);
  not NOT_2128(WX6370,WX6177);
  not NOT_2129(WX6372,WX6371);
  not NOT_2130(WX6373,WX6372);
  not NOT_2131(WX6377,WX6177);
  not NOT_2132(WX6379,WX6378);
  not NOT_2133(WX6380,WX6379);
  not NOT_2134(WX6384,WX6177);
  not NOT_2135(WX6386,WX6385);
  not NOT_2136(WX6387,WX6386);
  not NOT_2137(WX6391,WX6177);
  not NOT_2138(WX6393,WX6392);
  not NOT_2139(WX6394,WX6393);
  not NOT_2140(WX6398,WX6177);
  not NOT_2141(WX6400,WX6399);
  not NOT_2142(WX6401,WX6400);
  not NOT_2143(WX6402,RESET);
  not NOT_2144(WX6435,WX6402);
  not NOT_2145(WX6502,WX7468);
  not NOT_2146(WX6506,WX7469);
  not NOT_2147(WX6510,WX7469);
  not NOT_2148(WX6512,WX6503);
  not NOT_2149(WX6513,WX6512);
  not NOT_2150(WX6516,WX7468);
  not NOT_2151(WX6520,WX7469);
  not NOT_2152(WX6524,WX7469);
  not NOT_2153(WX6526,WX6517);
  not NOT_2154(WX6527,WX6526);
  not NOT_2155(WX6530,WX7468);
  not NOT_2156(WX6534,WX7469);
  not NOT_2157(WX6538,WX7469);
  not NOT_2158(WX6540,WX6531);
  not NOT_2159(WX6541,WX6540);
  not NOT_2160(WX6544,WX7468);
  not NOT_2161(WX6548,WX7469);
  not NOT_2162(WX6552,WX7469);
  not NOT_2163(WX6554,WX6545);
  not NOT_2164(WX6555,WX6554);
  not NOT_2165(WX6558,WX7468);
  not NOT_2166(WX6562,WX7469);
  not NOT_2167(WX6566,WX7469);
  not NOT_2168(WX6568,WX6559);
  not NOT_2169(WX6569,WX6568);
  not NOT_2170(WX6572,WX7468);
  not NOT_2171(WX6576,WX7469);
  not NOT_2172(WX6580,WX7469);
  not NOT_2173(WX6582,WX6573);
  not NOT_2174(WX6583,WX6582);
  not NOT_2175(WX6586,WX7468);
  not NOT_2176(WX6590,WX7469);
  not NOT_2177(WX6594,WX7469);
  not NOT_2178(WX6596,WX6587);
  not NOT_2179(WX6597,WX6596);
  not NOT_2180(WX6600,WX7468);
  not NOT_2181(WX6604,WX7469);
  not NOT_2182(WX6608,WX7469);
  not NOT_2183(WX6610,WX6601);
  not NOT_2184(WX6611,WX6610);
  not NOT_2185(WX6614,WX7468);
  not NOT_2186(WX6618,WX7469);
  not NOT_2187(WX6622,WX7469);
  not NOT_2188(WX6624,WX6615);
  not NOT_2189(WX6625,WX6624);
  not NOT_2190(WX6628,WX7468);
  not NOT_2191(WX6632,WX7469);
  not NOT_2192(WX6636,WX7469);
  not NOT_2193(WX6638,WX6629);
  not NOT_2194(WX6639,WX6638);
  not NOT_2195(WX6642,WX7468);
  not NOT_2196(WX6646,WX7469);
  not NOT_2197(WX6650,WX7469);
  not NOT_2198(WX6652,WX6643);
  not NOT_2199(WX6653,WX6652);
  not NOT_2200(WX6656,WX7468);
  not NOT_2201(WX6660,WX7469);
  not NOT_2202(WX6664,WX7469);
  not NOT_2203(WX6666,WX6657);
  not NOT_2204(WX6667,WX6666);
  not NOT_2205(WX6670,WX7468);
  not NOT_2206(WX6674,WX7469);
  not NOT_2207(WX6678,WX7469);
  not NOT_2208(WX6680,WX6671);
  not NOT_2209(WX6681,WX6680);
  not NOT_2210(WX6684,WX7468);
  not NOT_2211(WX6688,WX7469);
  not NOT_2212(WX6692,WX7469);
  not NOT_2213(WX6694,WX6685);
  not NOT_2214(WX6695,WX6694);
  not NOT_2215(WX6698,WX7468);
  not NOT_2216(WX6702,WX7469);
  not NOT_2217(WX6706,WX7469);
  not NOT_2218(WX6708,WX6699);
  not NOT_2219(WX6709,WX6708);
  not NOT_2220(WX6712,WX7468);
  not NOT_2221(WX6716,WX7469);
  not NOT_2222(WX6720,WX7469);
  not NOT_2223(WX6722,WX6713);
  not NOT_2224(WX6723,WX6722);
  not NOT_2225(WX6726,WX7468);
  not NOT_2226(WX6730,WX7469);
  not NOT_2227(WX6734,WX7469);
  not NOT_2228(WX6736,WX6727);
  not NOT_2229(WX6737,WX6736);
  not NOT_2230(WX6740,WX7468);
  not NOT_2231(WX6744,WX7469);
  not NOT_2232(WX6748,WX7469);
  not NOT_2233(WX6750,WX6741);
  not NOT_2234(WX6751,WX6750);
  not NOT_2235(WX6754,WX7468);
  not NOT_2236(WX6758,WX7469);
  not NOT_2237(WX6762,WX7469);
  not NOT_2238(WX6764,WX6755);
  not NOT_2239(WX6765,WX6764);
  not NOT_2240(WX6768,WX7468);
  not NOT_2241(WX6772,WX7469);
  not NOT_2242(WX6776,WX7469);
  not NOT_2243(WX6778,WX6769);
  not NOT_2244(WX6779,WX6778);
  not NOT_2245(WX6782,WX7468);
  not NOT_2246(WX6786,WX7469);
  not NOT_2247(WX6790,WX7469);
  not NOT_2248(WX6792,WX6783);
  not NOT_2249(WX6793,WX6792);
  not NOT_2250(WX6796,WX7468);
  not NOT_2251(WX6800,WX7469);
  not NOT_2252(WX6804,WX7469);
  not NOT_2253(WX6806,WX6797);
  not NOT_2254(WX6807,WX6806);
  not NOT_2255(WX6810,WX7468);
  not NOT_2256(WX6814,WX7469);
  not NOT_2257(WX6818,WX7469);
  not NOT_2258(WX6820,WX6811);
  not NOT_2259(WX6821,WX6820);
  not NOT_2260(WX6824,WX7468);
  not NOT_2261(WX6828,WX7469);
  not NOT_2262(WX6832,WX7469);
  not NOT_2263(WX6834,WX6825);
  not NOT_2264(WX6835,WX6834);
  not NOT_2265(WX6838,WX7468);
  not NOT_2266(WX6842,WX7469);
  not NOT_2267(WX6846,WX7469);
  not NOT_2268(WX6848,WX6839);
  not NOT_2269(WX6849,WX6848);
  not NOT_2270(WX6852,WX7468);
  not NOT_2271(WX6856,WX7469);
  not NOT_2272(WX6860,WX7469);
  not NOT_2273(WX6862,WX6853);
  not NOT_2274(WX6863,WX6862);
  not NOT_2275(WX6866,WX7468);
  not NOT_2276(WX6870,WX7469);
  not NOT_2277(WX6874,WX7469);
  not NOT_2278(WX6876,WX6867);
  not NOT_2279(WX6877,WX6876);
  not NOT_2280(WX6880,WX7468);
  not NOT_2281(WX6884,WX7469);
  not NOT_2282(WX6888,WX7469);
  not NOT_2283(WX6890,WX6881);
  not NOT_2284(WX6891,WX6890);
  not NOT_2285(WX6894,WX7468);
  not NOT_2286(WX6898,WX7469);
  not NOT_2287(WX6902,WX7469);
  not NOT_2288(WX6904,WX6895);
  not NOT_2289(WX6905,WX6904);
  not NOT_2290(WX6908,WX7468);
  not NOT_2291(WX6912,WX7469);
  not NOT_2292(WX6916,WX7469);
  not NOT_2293(WX6918,WX6909);
  not NOT_2294(WX6919,WX6918);
  not NOT_2295(WX6922,WX7468);
  not NOT_2296(WX6926,WX7469);
  not NOT_2297(WX6930,WX7469);
  not NOT_2298(WX6932,WX6923);
  not NOT_2299(WX6933,WX6932);
  not NOT_2300(WX6936,WX7468);
  not NOT_2301(WX6940,WX7469);
  not NOT_2302(WX6944,WX7469);
  not NOT_2303(WX6946,WX6937);
  not NOT_2304(WX6947,WX6946);
  not NOT_2305(WX6948,WX6950);
  not NOT_2306(WX7013,WX7430);
  not NOT_2307(WX7014,WX7432);
  not NOT_2308(WX7015,WX7434);
  not NOT_2309(WX7016,WX7436);
  not NOT_2310(WX7017,WX7438);
  not NOT_2311(WX7018,WX7440);
  not NOT_2312(WX7019,WX7442);
  not NOT_2313(WX7020,WX7444);
  not NOT_2314(WX7021,WX7446);
  not NOT_2315(WX7022,WX7448);
  not NOT_2316(WX7023,WX7450);
  not NOT_2317(WX7024,WX7452);
  not NOT_2318(WX7025,WX7454);
  not NOT_2319(WX7026,WX7456);
  not NOT_2320(WX7027,WX7458);
  not NOT_2321(WX7028,WX7460);
  not NOT_2322(WX7029,WX7398);
  not NOT_2323(WX7030,WX7400);
  not NOT_2324(WX7031,WX7402);
  not NOT_2325(WX7032,WX7404);
  not NOT_2326(WX7033,WX7406);
  not NOT_2327(WX7034,WX7408);
  not NOT_2328(WX7035,WX7410);
  not NOT_2329(WX7036,WX7412);
  not NOT_2330(WX7037,WX7414);
  not NOT_2331(WX7038,WX7416);
  not NOT_2332(WX7039,WX7418);
  not NOT_2333(WX7040,WX7420);
  not NOT_2334(WX7041,WX7422);
  not NOT_2335(WX7042,WX7424);
  not NOT_2336(WX7043,WX7426);
  not NOT_2337(WX7044,WX7428);
  not NOT_2338(WX7045,WX7013);
  not NOT_2339(WX7046,WX7014);
  not NOT_2340(WX7047,WX7015);
  not NOT_2341(WX7048,WX7016);
  not NOT_2342(WX7049,WX7017);
  not NOT_2343(WX7050,WX7018);
  not NOT_2344(WX7051,WX7019);
  not NOT_2345(WX7052,WX7020);
  not NOT_2346(WX7053,WX7021);
  not NOT_2347(WX7054,WX7022);
  not NOT_2348(WX7055,WX7023);
  not NOT_2349(WX7056,WX7024);
  not NOT_2350(WX7057,WX7025);
  not NOT_2351(WX7058,WX7026);
  not NOT_2352(WX7059,WX7027);
  not NOT_2353(WX7060,WX7028);
  not NOT_2354(WX7061,WX7029);
  not NOT_2355(WX7062,WX7030);
  not NOT_2356(WX7063,WX7031);
  not NOT_2357(WX7064,WX7032);
  not NOT_2358(WX7065,WX7033);
  not NOT_2359(WX7066,WX7034);
  not NOT_2360(WX7067,WX7035);
  not NOT_2361(WX7068,WX7036);
  not NOT_2362(WX7069,WX7037);
  not NOT_2363(WX7070,WX7038);
  not NOT_2364(WX7071,WX7039);
  not NOT_2365(WX7072,WX7040);
  not NOT_2366(WX7073,WX7041);
  not NOT_2367(WX7074,WX7042);
  not NOT_2368(WX7075,WX7043);
  not NOT_2369(WX7076,WX7044);
  not NOT_2370(WX7077,WX7302);
  not NOT_2371(WX7078,WX7304);
  not NOT_2372(WX7079,WX7306);
  not NOT_2373(WX7080,WX7308);
  not NOT_2374(WX7081,WX7310);
  not NOT_2375(WX7082,WX7312);
  not NOT_2376(WX7083,WX7314);
  not NOT_2377(WX7084,WX7316);
  not NOT_2378(WX7085,WX7318);
  not NOT_2379(WX7086,WX7320);
  not NOT_2380(WX7087,WX7322);
  not NOT_2381(WX7088,WX7324);
  not NOT_2382(WX7089,WX7326);
  not NOT_2383(WX7090,WX7328);
  not NOT_2384(WX7091,WX7330);
  not NOT_2385(WX7092,WX7332);
  not NOT_2386(WX7093,WX7334);
  not NOT_2387(WX7094,WX7336);
  not NOT_2388(WX7095,WX7338);
  not NOT_2389(WX7096,WX7340);
  not NOT_2390(WX7097,WX7342);
  not NOT_2391(WX7098,WX7344);
  not NOT_2392(WX7099,WX7346);
  not NOT_2393(WX7100,WX7348);
  not NOT_2394(WX7101,WX7350);
  not NOT_2395(WX7102,WX7352);
  not NOT_2396(WX7103,WX7354);
  not NOT_2397(WX7104,WX7356);
  not NOT_2398(WX7105,WX7358);
  not NOT_2399(WX7106,WX7360);
  not NOT_2400(WX7107,WX7362);
  not NOT_2401(WX7108,WX7364);
  not NOT_2402(WX7397,WX7381);
  not NOT_2403(WX7398,WX7397);
  not NOT_2404(WX7399,WX7382);
  not NOT_2405(WX7400,WX7399);
  not NOT_2406(WX7401,WX7383);
  not NOT_2407(WX7402,WX7401);
  not NOT_2408(WX7403,WX7384);
  not NOT_2409(WX7404,WX7403);
  not NOT_2410(WX7405,WX7385);
  not NOT_2411(WX7406,WX7405);
  not NOT_2412(WX7407,WX7386);
  not NOT_2413(WX7408,WX7407);
  not NOT_2414(WX7409,WX7387);
  not NOT_2415(WX7410,WX7409);
  not NOT_2416(WX7411,WX7388);
  not NOT_2417(WX7412,WX7411);
  not NOT_2418(WX7413,WX7389);
  not NOT_2419(WX7414,WX7413);
  not NOT_2420(WX7415,WX7390);
  not NOT_2421(WX7416,WX7415);
  not NOT_2422(WX7417,WX7391);
  not NOT_2423(WX7418,WX7417);
  not NOT_2424(WX7419,WX7392);
  not NOT_2425(WX7420,WX7419);
  not NOT_2426(WX7421,WX7393);
  not NOT_2427(WX7422,WX7421);
  not NOT_2428(WX7423,WX7394);
  not NOT_2429(WX7424,WX7423);
  not NOT_2430(WX7425,WX7395);
  not NOT_2431(WX7426,WX7425);
  not NOT_2432(WX7427,WX7396);
  not NOT_2433(WX7428,WX7427);
  not NOT_2434(WX7429,WX7365);
  not NOT_2435(WX7430,WX7429);
  not NOT_2436(WX7431,WX7366);
  not NOT_2437(WX7432,WX7431);
  not NOT_2438(WX7433,WX7367);
  not NOT_2439(WX7434,WX7433);
  not NOT_2440(WX7435,WX7368);
  not NOT_2441(WX7436,WX7435);
  not NOT_2442(WX7437,WX7369);
  not NOT_2443(WX7438,WX7437);
  not NOT_2444(WX7439,WX7370);
  not NOT_2445(WX7440,WX7439);
  not NOT_2446(WX7441,WX7371);
  not NOT_2447(WX7442,WX7441);
  not NOT_2448(WX7443,WX7372);
  not NOT_2449(WX7444,WX7443);
  not NOT_2450(WX7445,WX7373);
  not NOT_2451(WX7446,WX7445);
  not NOT_2452(WX7447,WX7374);
  not NOT_2453(WX7448,WX7447);
  not NOT_2454(WX7449,WX7375);
  not NOT_2455(WX7450,WX7449);
  not NOT_2456(WX7451,WX7376);
  not NOT_2457(WX7452,WX7451);
  not NOT_2458(WX7453,WX7377);
  not NOT_2459(WX7454,WX7453);
  not NOT_2460(WX7455,WX7378);
  not NOT_2461(WX7456,WX7455);
  not NOT_2462(WX7457,WX7379);
  not NOT_2463(WX7458,WX7457);
  not NOT_2464(WX7459,WX7380);
  not NOT_2465(WX7460,WX7459);
  not NOT_2466(WX7461,TM0);
  not NOT_2467(WX7462,TM0);
  not NOT_2468(WX7463,TM0);
  not NOT_2469(WX7464,TM1);
  not NOT_2470(WX7465,TM1);
  not NOT_2471(WX7466,WX7465);
  not NOT_2472(WX7467,WX7463);
  not NOT_2473(WX7468,WX7464);
  not NOT_2474(WX7469,WX7462);
  not NOT_2475(WX7470,WX7461);
  not NOT_2476(WX7474,WX7470);
  not NOT_2477(WX7476,WX7475);
  not NOT_2478(WX7477,WX7476);
  not NOT_2479(WX7481,WX7470);
  not NOT_2480(WX7483,WX7482);
  not NOT_2481(WX7484,WX7483);
  not NOT_2482(WX7488,WX7470);
  not NOT_2483(WX7490,WX7489);
  not NOT_2484(WX7491,WX7490);
  not NOT_2485(WX7495,WX7470);
  not NOT_2486(WX7497,WX7496);
  not NOT_2487(WX7498,WX7497);
  not NOT_2488(WX7502,WX7470);
  not NOT_2489(WX7504,WX7503);
  not NOT_2490(WX7505,WX7504);
  not NOT_2491(WX7509,WX7470);
  not NOT_2492(WX7511,WX7510);
  not NOT_2493(WX7512,WX7511);
  not NOT_2494(WX7516,WX7470);
  not NOT_2495(WX7518,WX7517);
  not NOT_2496(WX7519,WX7518);
  not NOT_2497(WX7523,WX7470);
  not NOT_2498(WX7525,WX7524);
  not NOT_2499(WX7526,WX7525);
  not NOT_2500(WX7530,WX7470);
  not NOT_2501(WX7532,WX7531);
  not NOT_2502(WX7533,WX7532);
  not NOT_2503(WX7537,WX7470);
  not NOT_2504(WX7539,WX7538);
  not NOT_2505(WX7540,WX7539);
  not NOT_2506(WX7544,WX7470);
  not NOT_2507(WX7546,WX7545);
  not NOT_2508(WX7547,WX7546);
  not NOT_2509(WX7551,WX7470);
  not NOT_2510(WX7553,WX7552);
  not NOT_2511(WX7554,WX7553);
  not NOT_2512(WX7558,WX7470);
  not NOT_2513(WX7560,WX7559);
  not NOT_2514(WX7561,WX7560);
  not NOT_2515(WX7565,WX7470);
  not NOT_2516(WX7567,WX7566);
  not NOT_2517(WX7568,WX7567);
  not NOT_2518(WX7572,WX7470);
  not NOT_2519(WX7574,WX7573);
  not NOT_2520(WX7575,WX7574);
  not NOT_2521(WX7579,WX7470);
  not NOT_2522(WX7581,WX7580);
  not NOT_2523(WX7582,WX7581);
  not NOT_2524(WX7586,WX7470);
  not NOT_2525(WX7588,WX7587);
  not NOT_2526(WX7589,WX7588);
  not NOT_2527(WX7593,WX7470);
  not NOT_2528(WX7595,WX7594);
  not NOT_2529(WX7596,WX7595);
  not NOT_2530(WX7600,WX7470);
  not NOT_2531(WX7602,WX7601);
  not NOT_2532(WX7603,WX7602);
  not NOT_2533(WX7607,WX7470);
  not NOT_2534(WX7609,WX7608);
  not NOT_2535(WX7610,WX7609);
  not NOT_2536(WX7614,WX7470);
  not NOT_2537(WX7616,WX7615);
  not NOT_2538(WX7617,WX7616);
  not NOT_2539(WX7621,WX7470);
  not NOT_2540(WX7623,WX7622);
  not NOT_2541(WX7624,WX7623);
  not NOT_2542(WX7628,WX7470);
  not NOT_2543(WX7630,WX7629);
  not NOT_2544(WX7631,WX7630);
  not NOT_2545(WX7635,WX7470);
  not NOT_2546(WX7637,WX7636);
  not NOT_2547(WX7638,WX7637);
  not NOT_2548(WX7642,WX7470);
  not NOT_2549(WX7644,WX7643);
  not NOT_2550(WX7645,WX7644);
  not NOT_2551(WX7649,WX7470);
  not NOT_2552(WX7651,WX7650);
  not NOT_2553(WX7652,WX7651);
  not NOT_2554(WX7656,WX7470);
  not NOT_2555(WX7658,WX7657);
  not NOT_2556(WX7659,WX7658);
  not NOT_2557(WX7663,WX7470);
  not NOT_2558(WX7665,WX7664);
  not NOT_2559(WX7666,WX7665);
  not NOT_2560(WX7670,WX7470);
  not NOT_2561(WX7672,WX7671);
  not NOT_2562(WX7673,WX7672);
  not NOT_2563(WX7677,WX7470);
  not NOT_2564(WX7679,WX7678);
  not NOT_2565(WX7680,WX7679);
  not NOT_2566(WX7684,WX7470);
  not NOT_2567(WX7686,WX7685);
  not NOT_2568(WX7687,WX7686);
  not NOT_2569(WX7691,WX7470);
  not NOT_2570(WX7693,WX7692);
  not NOT_2571(WX7694,WX7693);
  not NOT_2572(WX7695,RESET);
  not NOT_2573(WX7728,WX7695);
  not NOT_2574(WX7795,WX8761);
  not NOT_2575(WX7799,WX8762);
  not NOT_2576(WX7803,WX8762);
  not NOT_2577(WX7805,WX7796);
  not NOT_2578(WX7806,WX7805);
  not NOT_2579(WX7809,WX8761);
  not NOT_2580(WX7813,WX8762);
  not NOT_2581(WX7817,WX8762);
  not NOT_2582(WX7819,WX7810);
  not NOT_2583(WX7820,WX7819);
  not NOT_2584(WX7823,WX8761);
  not NOT_2585(WX7827,WX8762);
  not NOT_2586(WX7831,WX8762);
  not NOT_2587(WX7833,WX7824);
  not NOT_2588(WX7834,WX7833);
  not NOT_2589(WX7837,WX8761);
  not NOT_2590(WX7841,WX8762);
  not NOT_2591(WX7845,WX8762);
  not NOT_2592(WX7847,WX7838);
  not NOT_2593(WX7848,WX7847);
  not NOT_2594(WX7851,WX8761);
  not NOT_2595(WX7855,WX8762);
  not NOT_2596(WX7859,WX8762);
  not NOT_2597(WX7861,WX7852);
  not NOT_2598(WX7862,WX7861);
  not NOT_2599(WX7865,WX8761);
  not NOT_2600(WX7869,WX8762);
  not NOT_2601(WX7873,WX8762);
  not NOT_2602(WX7875,WX7866);
  not NOT_2603(WX7876,WX7875);
  not NOT_2604(WX7879,WX8761);
  not NOT_2605(WX7883,WX8762);
  not NOT_2606(WX7887,WX8762);
  not NOT_2607(WX7889,WX7880);
  not NOT_2608(WX7890,WX7889);
  not NOT_2609(WX7893,WX8761);
  not NOT_2610(WX7897,WX8762);
  not NOT_2611(WX7901,WX8762);
  not NOT_2612(WX7903,WX7894);
  not NOT_2613(WX7904,WX7903);
  not NOT_2614(WX7907,WX8761);
  not NOT_2615(WX7911,WX8762);
  not NOT_2616(WX7915,WX8762);
  not NOT_2617(WX7917,WX7908);
  not NOT_2618(WX7918,WX7917);
  not NOT_2619(WX7921,WX8761);
  not NOT_2620(WX7925,WX8762);
  not NOT_2621(WX7929,WX8762);
  not NOT_2622(WX7931,WX7922);
  not NOT_2623(WX7932,WX7931);
  not NOT_2624(WX7935,WX8761);
  not NOT_2625(WX7939,WX8762);
  not NOT_2626(WX7943,WX8762);
  not NOT_2627(WX7945,WX7936);
  not NOT_2628(WX7946,WX7945);
  not NOT_2629(WX7949,WX8761);
  not NOT_2630(WX7953,WX8762);
  not NOT_2631(WX7957,WX8762);
  not NOT_2632(WX7959,WX7950);
  not NOT_2633(WX7960,WX7959);
  not NOT_2634(WX7963,WX8761);
  not NOT_2635(WX7967,WX8762);
  not NOT_2636(WX7971,WX8762);
  not NOT_2637(WX7973,WX7964);
  not NOT_2638(WX7974,WX7973);
  not NOT_2639(WX7977,WX8761);
  not NOT_2640(WX7981,WX8762);
  not NOT_2641(WX7985,WX8762);
  not NOT_2642(WX7987,WX7978);
  not NOT_2643(WX7988,WX7987);
  not NOT_2644(WX7991,WX8761);
  not NOT_2645(WX7995,WX8762);
  not NOT_2646(WX7999,WX8762);
  not NOT_2647(WX8001,WX7992);
  not NOT_2648(WX8002,WX8001);
  not NOT_2649(WX8005,WX8761);
  not NOT_2650(WX8009,WX8762);
  not NOT_2651(WX8013,WX8762);
  not NOT_2652(WX8015,WX8006);
  not NOT_2653(WX8016,WX8015);
  not NOT_2654(WX8019,WX8761);
  not NOT_2655(WX8023,WX8762);
  not NOT_2656(WX8027,WX8762);
  not NOT_2657(WX8029,WX8020);
  not NOT_2658(WX8030,WX8029);
  not NOT_2659(WX8033,WX8761);
  not NOT_2660(WX8037,WX8762);
  not NOT_2661(WX8041,WX8762);
  not NOT_2662(WX8043,WX8034);
  not NOT_2663(WX8044,WX8043);
  not NOT_2664(WX8047,WX8761);
  not NOT_2665(WX8051,WX8762);
  not NOT_2666(WX8055,WX8762);
  not NOT_2667(WX8057,WX8048);
  not NOT_2668(WX8058,WX8057);
  not NOT_2669(WX8061,WX8761);
  not NOT_2670(WX8065,WX8762);
  not NOT_2671(WX8069,WX8762);
  not NOT_2672(WX8071,WX8062);
  not NOT_2673(WX8072,WX8071);
  not NOT_2674(WX8075,WX8761);
  not NOT_2675(WX8079,WX8762);
  not NOT_2676(WX8083,WX8762);
  not NOT_2677(WX8085,WX8076);
  not NOT_2678(WX8086,WX8085);
  not NOT_2679(WX8089,WX8761);
  not NOT_2680(WX8093,WX8762);
  not NOT_2681(WX8097,WX8762);
  not NOT_2682(WX8099,WX8090);
  not NOT_2683(WX8100,WX8099);
  not NOT_2684(WX8103,WX8761);
  not NOT_2685(WX8107,WX8762);
  not NOT_2686(WX8111,WX8762);
  not NOT_2687(WX8113,WX8104);
  not NOT_2688(WX8114,WX8113);
  not NOT_2689(WX8117,WX8761);
  not NOT_2690(WX8121,WX8762);
  not NOT_2691(WX8125,WX8762);
  not NOT_2692(WX8127,WX8118);
  not NOT_2693(WX8128,WX8127);
  not NOT_2694(WX8131,WX8761);
  not NOT_2695(WX8135,WX8762);
  not NOT_2696(WX8139,WX8762);
  not NOT_2697(WX8141,WX8132);
  not NOT_2698(WX8142,WX8141);
  not NOT_2699(WX8145,WX8761);
  not NOT_2700(WX8149,WX8762);
  not NOT_2701(WX8153,WX8762);
  not NOT_2702(WX8155,WX8146);
  not NOT_2703(WX8156,WX8155);
  not NOT_2704(WX8159,WX8761);
  not NOT_2705(WX8163,WX8762);
  not NOT_2706(WX8167,WX8762);
  not NOT_2707(WX8169,WX8160);
  not NOT_2708(WX8170,WX8169);
  not NOT_2709(WX8173,WX8761);
  not NOT_2710(WX8177,WX8762);
  not NOT_2711(WX8181,WX8762);
  not NOT_2712(WX8183,WX8174);
  not NOT_2713(WX8184,WX8183);
  not NOT_2714(WX8187,WX8761);
  not NOT_2715(WX8191,WX8762);
  not NOT_2716(WX8195,WX8762);
  not NOT_2717(WX8197,WX8188);
  not NOT_2718(WX8198,WX8197);
  not NOT_2719(WX8201,WX8761);
  not NOT_2720(WX8205,WX8762);
  not NOT_2721(WX8209,WX8762);
  not NOT_2722(WX8211,WX8202);
  not NOT_2723(WX8212,WX8211);
  not NOT_2724(WX8215,WX8761);
  not NOT_2725(WX8219,WX8762);
  not NOT_2726(WX8223,WX8762);
  not NOT_2727(WX8225,WX8216);
  not NOT_2728(WX8226,WX8225);
  not NOT_2729(WX8229,WX8761);
  not NOT_2730(WX8233,WX8762);
  not NOT_2731(WX8237,WX8762);
  not NOT_2732(WX8239,WX8230);
  not NOT_2733(WX8240,WX8239);
  not NOT_2734(WX8241,WX8243);
  not NOT_2735(WX8306,WX8723);
  not NOT_2736(WX8307,WX8725);
  not NOT_2737(WX8308,WX8727);
  not NOT_2738(WX8309,WX8729);
  not NOT_2739(WX8310,WX8731);
  not NOT_2740(WX8311,WX8733);
  not NOT_2741(WX8312,WX8735);
  not NOT_2742(WX8313,WX8737);
  not NOT_2743(WX8314,WX8739);
  not NOT_2744(WX8315,WX8741);
  not NOT_2745(WX8316,WX8743);
  not NOT_2746(WX8317,WX8745);
  not NOT_2747(WX8318,WX8747);
  not NOT_2748(WX8319,WX8749);
  not NOT_2749(WX8320,WX8751);
  not NOT_2750(WX8321,WX8753);
  not NOT_2751(WX8322,WX8691);
  not NOT_2752(WX8323,WX8693);
  not NOT_2753(WX8324,WX8695);
  not NOT_2754(WX8325,WX8697);
  not NOT_2755(WX8326,WX8699);
  not NOT_2756(WX8327,WX8701);
  not NOT_2757(WX8328,WX8703);
  not NOT_2758(WX8329,WX8705);
  not NOT_2759(WX8330,WX8707);
  not NOT_2760(WX8331,WX8709);
  not NOT_2761(WX8332,WX8711);
  not NOT_2762(WX8333,WX8713);
  not NOT_2763(WX8334,WX8715);
  not NOT_2764(WX8335,WX8717);
  not NOT_2765(WX8336,WX8719);
  not NOT_2766(WX8337,WX8721);
  not NOT_2767(WX8338,WX8306);
  not NOT_2768(WX8339,WX8307);
  not NOT_2769(WX8340,WX8308);
  not NOT_2770(WX8341,WX8309);
  not NOT_2771(WX8342,WX8310);
  not NOT_2772(WX8343,WX8311);
  not NOT_2773(WX8344,WX8312);
  not NOT_2774(WX8345,WX8313);
  not NOT_2775(WX8346,WX8314);
  not NOT_2776(WX8347,WX8315);
  not NOT_2777(WX8348,WX8316);
  not NOT_2778(WX8349,WX8317);
  not NOT_2779(WX8350,WX8318);
  not NOT_2780(WX8351,WX8319);
  not NOT_2781(WX8352,WX8320);
  not NOT_2782(WX8353,WX8321);
  not NOT_2783(WX8354,WX8322);
  not NOT_2784(WX8355,WX8323);
  not NOT_2785(WX8356,WX8324);
  not NOT_2786(WX8357,WX8325);
  not NOT_2787(WX8358,WX8326);
  not NOT_2788(WX8359,WX8327);
  not NOT_2789(WX8360,WX8328);
  not NOT_2790(WX8361,WX8329);
  not NOT_2791(WX8362,WX8330);
  not NOT_2792(WX8363,WX8331);
  not NOT_2793(WX8364,WX8332);
  not NOT_2794(WX8365,WX8333);
  not NOT_2795(WX8366,WX8334);
  not NOT_2796(WX8367,WX8335);
  not NOT_2797(WX8368,WX8336);
  not NOT_2798(WX8369,WX8337);
  not NOT_2799(WX8370,WX8595);
  not NOT_2800(WX8371,WX8597);
  not NOT_2801(WX8372,WX8599);
  not NOT_2802(WX8373,WX8601);
  not NOT_2803(WX8374,WX8603);
  not NOT_2804(WX8375,WX8605);
  not NOT_2805(WX8376,WX8607);
  not NOT_2806(WX8377,WX8609);
  not NOT_2807(WX8378,WX8611);
  not NOT_2808(WX8379,WX8613);
  not NOT_2809(WX8380,WX8615);
  not NOT_2810(WX8381,WX8617);
  not NOT_2811(WX8382,WX8619);
  not NOT_2812(WX8383,WX8621);
  not NOT_2813(WX8384,WX8623);
  not NOT_2814(WX8385,WX8625);
  not NOT_2815(WX8386,WX8627);
  not NOT_2816(WX8387,WX8629);
  not NOT_2817(WX8388,WX8631);
  not NOT_2818(WX8389,WX8633);
  not NOT_2819(WX8390,WX8635);
  not NOT_2820(WX8391,WX8637);
  not NOT_2821(WX8392,WX8639);
  not NOT_2822(WX8393,WX8641);
  not NOT_2823(WX8394,WX8643);
  not NOT_2824(WX8395,WX8645);
  not NOT_2825(WX8396,WX8647);
  not NOT_2826(WX8397,WX8649);
  not NOT_2827(WX8398,WX8651);
  not NOT_2828(WX8399,WX8653);
  not NOT_2829(WX8400,WX8655);
  not NOT_2830(WX8401,WX8657);
  not NOT_2831(WX8690,WX8674);
  not NOT_2832(WX8691,WX8690);
  not NOT_2833(WX8692,WX8675);
  not NOT_2834(WX8693,WX8692);
  not NOT_2835(WX8694,WX8676);
  not NOT_2836(WX8695,WX8694);
  not NOT_2837(WX8696,WX8677);
  not NOT_2838(WX8697,WX8696);
  not NOT_2839(WX8698,WX8678);
  not NOT_2840(WX8699,WX8698);
  not NOT_2841(WX8700,WX8679);
  not NOT_2842(WX8701,WX8700);
  not NOT_2843(WX8702,WX8680);
  not NOT_2844(WX8703,WX8702);
  not NOT_2845(WX8704,WX8681);
  not NOT_2846(WX8705,WX8704);
  not NOT_2847(WX8706,WX8682);
  not NOT_2848(WX8707,WX8706);
  not NOT_2849(WX8708,WX8683);
  not NOT_2850(WX8709,WX8708);
  not NOT_2851(WX8710,WX8684);
  not NOT_2852(WX8711,WX8710);
  not NOT_2853(WX8712,WX8685);
  not NOT_2854(WX8713,WX8712);
  not NOT_2855(WX8714,WX8686);
  not NOT_2856(WX8715,WX8714);
  not NOT_2857(WX8716,WX8687);
  not NOT_2858(WX8717,WX8716);
  not NOT_2859(WX8718,WX8688);
  not NOT_2860(WX8719,WX8718);
  not NOT_2861(WX8720,WX8689);
  not NOT_2862(WX8721,WX8720);
  not NOT_2863(WX8722,WX8658);
  not NOT_2864(WX8723,WX8722);
  not NOT_2865(WX8724,WX8659);
  not NOT_2866(WX8725,WX8724);
  not NOT_2867(WX8726,WX8660);
  not NOT_2868(WX8727,WX8726);
  not NOT_2869(WX8728,WX8661);
  not NOT_2870(WX8729,WX8728);
  not NOT_2871(WX8730,WX8662);
  not NOT_2872(WX8731,WX8730);
  not NOT_2873(WX8732,WX8663);
  not NOT_2874(WX8733,WX8732);
  not NOT_2875(WX8734,WX8664);
  not NOT_2876(WX8735,WX8734);
  not NOT_2877(WX8736,WX8665);
  not NOT_2878(WX8737,WX8736);
  not NOT_2879(WX8738,WX8666);
  not NOT_2880(WX8739,WX8738);
  not NOT_2881(WX8740,WX8667);
  not NOT_2882(WX8741,WX8740);
  not NOT_2883(WX8742,WX8668);
  not NOT_2884(WX8743,WX8742);
  not NOT_2885(WX8744,WX8669);
  not NOT_2886(WX8745,WX8744);
  not NOT_2887(WX8746,WX8670);
  not NOT_2888(WX8747,WX8746);
  not NOT_2889(WX8748,WX8671);
  not NOT_2890(WX8749,WX8748);
  not NOT_2891(WX8750,WX8672);
  not NOT_2892(WX8751,WX8750);
  not NOT_2893(WX8752,WX8673);
  not NOT_2894(WX8753,WX8752);
  not NOT_2895(WX8754,TM0);
  not NOT_2896(WX8755,TM0);
  not NOT_2897(WX8756,TM0);
  not NOT_2898(WX8757,TM1);
  not NOT_2899(WX8758,TM1);
  not NOT_2900(WX8759,WX8758);
  not NOT_2901(WX8760,WX8756);
  not NOT_2902(WX8761,WX8757);
  not NOT_2903(WX8762,WX8755);
  not NOT_2904(WX8763,WX8754);
  not NOT_2905(WX8767,WX8763);
  not NOT_2906(WX8769,WX8768);
  not NOT_2907(WX8770,WX8769);
  not NOT_2908(WX8774,WX8763);
  not NOT_2909(WX8776,WX8775);
  not NOT_2910(WX8777,WX8776);
  not NOT_2911(WX8781,WX8763);
  not NOT_2912(WX8783,WX8782);
  not NOT_2913(WX8784,WX8783);
  not NOT_2914(WX8788,WX8763);
  not NOT_2915(WX8790,WX8789);
  not NOT_2916(WX8791,WX8790);
  not NOT_2917(WX8795,WX8763);
  not NOT_2918(WX8797,WX8796);
  not NOT_2919(WX8798,WX8797);
  not NOT_2920(WX8802,WX8763);
  not NOT_2921(WX8804,WX8803);
  not NOT_2922(WX8805,WX8804);
  not NOT_2923(WX8809,WX8763);
  not NOT_2924(WX8811,WX8810);
  not NOT_2925(WX8812,WX8811);
  not NOT_2926(WX8816,WX8763);
  not NOT_2927(WX8818,WX8817);
  not NOT_2928(WX8819,WX8818);
  not NOT_2929(WX8823,WX8763);
  not NOT_2930(WX8825,WX8824);
  not NOT_2931(WX8826,WX8825);
  not NOT_2932(WX8830,WX8763);
  not NOT_2933(WX8832,WX8831);
  not NOT_2934(WX8833,WX8832);
  not NOT_2935(WX8837,WX8763);
  not NOT_2936(WX8839,WX8838);
  not NOT_2937(WX8840,WX8839);
  not NOT_2938(WX8844,WX8763);
  not NOT_2939(WX8846,WX8845);
  not NOT_2940(WX8847,WX8846);
  not NOT_2941(WX8851,WX8763);
  not NOT_2942(WX8853,WX8852);
  not NOT_2943(WX8854,WX8853);
  not NOT_2944(WX8858,WX8763);
  not NOT_2945(WX8860,WX8859);
  not NOT_2946(WX8861,WX8860);
  not NOT_2947(WX8865,WX8763);
  not NOT_2948(WX8867,WX8866);
  not NOT_2949(WX8868,WX8867);
  not NOT_2950(WX8872,WX8763);
  not NOT_2951(WX8874,WX8873);
  not NOT_2952(WX8875,WX8874);
  not NOT_2953(WX8879,WX8763);
  not NOT_2954(WX8881,WX8880);
  not NOT_2955(WX8882,WX8881);
  not NOT_2956(WX8886,WX8763);
  not NOT_2957(WX8888,WX8887);
  not NOT_2958(WX8889,WX8888);
  not NOT_2959(WX8893,WX8763);
  not NOT_2960(WX8895,WX8894);
  not NOT_2961(WX8896,WX8895);
  not NOT_2962(WX8900,WX8763);
  not NOT_2963(WX8902,WX8901);
  not NOT_2964(WX8903,WX8902);
  not NOT_2965(WX8907,WX8763);
  not NOT_2966(WX8909,WX8908);
  not NOT_2967(WX8910,WX8909);
  not NOT_2968(WX8914,WX8763);
  not NOT_2969(WX8916,WX8915);
  not NOT_2970(WX8917,WX8916);
  not NOT_2971(WX8921,WX8763);
  not NOT_2972(WX8923,WX8922);
  not NOT_2973(WX8924,WX8923);
  not NOT_2974(WX8928,WX8763);
  not NOT_2975(WX8930,WX8929);
  not NOT_2976(WX8931,WX8930);
  not NOT_2977(WX8935,WX8763);
  not NOT_2978(WX8937,WX8936);
  not NOT_2979(WX8938,WX8937);
  not NOT_2980(WX8942,WX8763);
  not NOT_2981(WX8944,WX8943);
  not NOT_2982(WX8945,WX8944);
  not NOT_2983(WX8949,WX8763);
  not NOT_2984(WX8951,WX8950);
  not NOT_2985(WX8952,WX8951);
  not NOT_2986(WX8956,WX8763);
  not NOT_2987(WX8958,WX8957);
  not NOT_2988(WX8959,WX8958);
  not NOT_2989(WX8963,WX8763);
  not NOT_2990(WX8965,WX8964);
  not NOT_2991(WX8966,WX8965);
  not NOT_2992(WX8970,WX8763);
  not NOT_2993(WX8972,WX8971);
  not NOT_2994(WX8973,WX8972);
  not NOT_2995(WX8977,WX8763);
  not NOT_2996(WX8979,WX8978);
  not NOT_2997(WX8980,WX8979);
  not NOT_2998(WX8984,WX8763);
  not NOT_2999(WX8986,WX8985);
  not NOT_3000(WX8987,WX8986);
  not NOT_3001(WX8988,RESET);
  not NOT_3002(WX9021,WX8988);
  not NOT_3003(WX9088,WX10054);
  not NOT_3004(WX9092,WX10055);
  not NOT_3005(WX9096,WX10055);
  not NOT_3006(WX9098,WX9089);
  not NOT_3007(WX9099,WX9098);
  not NOT_3008(WX9102,WX10054);
  not NOT_3009(WX9106,WX10055);
  not NOT_3010(WX9110,WX10055);
  not NOT_3011(WX9112,WX9103);
  not NOT_3012(WX9113,WX9112);
  not NOT_3013(WX9116,WX10054);
  not NOT_3014(WX9120,WX10055);
  not NOT_3015(WX9124,WX10055);
  not NOT_3016(WX9126,WX9117);
  not NOT_3017(WX9127,WX9126);
  not NOT_3018(WX9130,WX10054);
  not NOT_3019(WX9134,WX10055);
  not NOT_3020(WX9138,WX10055);
  not NOT_3021(WX9140,WX9131);
  not NOT_3022(WX9141,WX9140);
  not NOT_3023(WX9144,WX10054);
  not NOT_3024(WX9148,WX10055);
  not NOT_3025(WX9152,WX10055);
  not NOT_3026(WX9154,WX9145);
  not NOT_3027(WX9155,WX9154);
  not NOT_3028(WX9158,WX10054);
  not NOT_3029(WX9162,WX10055);
  not NOT_3030(WX9166,WX10055);
  not NOT_3031(WX9168,WX9159);
  not NOT_3032(WX9169,WX9168);
  not NOT_3033(WX9172,WX10054);
  not NOT_3034(WX9176,WX10055);
  not NOT_3035(WX9180,WX10055);
  not NOT_3036(WX9182,WX9173);
  not NOT_3037(WX9183,WX9182);
  not NOT_3038(WX9186,WX10054);
  not NOT_3039(WX9190,WX10055);
  not NOT_3040(WX9194,WX10055);
  not NOT_3041(WX9196,WX9187);
  not NOT_3042(WX9197,WX9196);
  not NOT_3043(WX9200,WX10054);
  not NOT_3044(WX9204,WX10055);
  not NOT_3045(WX9208,WX10055);
  not NOT_3046(WX9210,WX9201);
  not NOT_3047(WX9211,WX9210);
  not NOT_3048(WX9214,WX10054);
  not NOT_3049(WX9218,WX10055);
  not NOT_3050(WX9222,WX10055);
  not NOT_3051(WX9224,WX9215);
  not NOT_3052(WX9225,WX9224);
  not NOT_3053(WX9228,WX10054);
  not NOT_3054(WX9232,WX10055);
  not NOT_3055(WX9236,WX10055);
  not NOT_3056(WX9238,WX9229);
  not NOT_3057(WX9239,WX9238);
  not NOT_3058(WX9242,WX10054);
  not NOT_3059(WX9246,WX10055);
  not NOT_3060(WX9250,WX10055);
  not NOT_3061(WX9252,WX9243);
  not NOT_3062(WX9253,WX9252);
  not NOT_3063(WX9256,WX10054);
  not NOT_3064(WX9260,WX10055);
  not NOT_3065(WX9264,WX10055);
  not NOT_3066(WX9266,WX9257);
  not NOT_3067(WX9267,WX9266);
  not NOT_3068(WX9270,WX10054);
  not NOT_3069(WX9274,WX10055);
  not NOT_3070(WX9278,WX10055);
  not NOT_3071(WX9280,WX9271);
  not NOT_3072(WX9281,WX9280);
  not NOT_3073(WX9284,WX10054);
  not NOT_3074(WX9288,WX10055);
  not NOT_3075(WX9292,WX10055);
  not NOT_3076(WX9294,WX9285);
  not NOT_3077(WX9295,WX9294);
  not NOT_3078(WX9298,WX10054);
  not NOT_3079(WX9302,WX10055);
  not NOT_3080(WX9306,WX10055);
  not NOT_3081(WX9308,WX9299);
  not NOT_3082(WX9309,WX9308);
  not NOT_3083(WX9312,WX10054);
  not NOT_3084(WX9316,WX10055);
  not NOT_3085(WX9320,WX10055);
  not NOT_3086(WX9322,WX9313);
  not NOT_3087(WX9323,WX9322);
  not NOT_3088(WX9326,WX10054);
  not NOT_3089(WX9330,WX10055);
  not NOT_3090(WX9334,WX10055);
  not NOT_3091(WX9336,WX9327);
  not NOT_3092(WX9337,WX9336);
  not NOT_3093(WX9340,WX10054);
  not NOT_3094(WX9344,WX10055);
  not NOT_3095(WX9348,WX10055);
  not NOT_3096(WX9350,WX9341);
  not NOT_3097(WX9351,WX9350);
  not NOT_3098(WX9354,WX10054);
  not NOT_3099(WX9358,WX10055);
  not NOT_3100(WX9362,WX10055);
  not NOT_3101(WX9364,WX9355);
  not NOT_3102(WX9365,WX9364);
  not NOT_3103(WX9368,WX10054);
  not NOT_3104(WX9372,WX10055);
  not NOT_3105(WX9376,WX10055);
  not NOT_3106(WX9378,WX9369);
  not NOT_3107(WX9379,WX9378);
  not NOT_3108(WX9382,WX10054);
  not NOT_3109(WX9386,WX10055);
  not NOT_3110(WX9390,WX10055);
  not NOT_3111(WX9392,WX9383);
  not NOT_3112(WX9393,WX9392);
  not NOT_3113(WX9396,WX10054);
  not NOT_3114(WX9400,WX10055);
  not NOT_3115(WX9404,WX10055);
  not NOT_3116(WX9406,WX9397);
  not NOT_3117(WX9407,WX9406);
  not NOT_3118(WX9410,WX10054);
  not NOT_3119(WX9414,WX10055);
  not NOT_3120(WX9418,WX10055);
  not NOT_3121(WX9420,WX9411);
  not NOT_3122(WX9421,WX9420);
  not NOT_3123(WX9424,WX10054);
  not NOT_3124(WX9428,WX10055);
  not NOT_3125(WX9432,WX10055);
  not NOT_3126(WX9434,WX9425);
  not NOT_3127(WX9435,WX9434);
  not NOT_3128(WX9438,WX10054);
  not NOT_3129(WX9442,WX10055);
  not NOT_3130(WX9446,WX10055);
  not NOT_3131(WX9448,WX9439);
  not NOT_3132(WX9449,WX9448);
  not NOT_3133(WX9452,WX10054);
  not NOT_3134(WX9456,WX10055);
  not NOT_3135(WX9460,WX10055);
  not NOT_3136(WX9462,WX9453);
  not NOT_3137(WX9463,WX9462);
  not NOT_3138(WX9466,WX10054);
  not NOT_3139(WX9470,WX10055);
  not NOT_3140(WX9474,WX10055);
  not NOT_3141(WX9476,WX9467);
  not NOT_3142(WX9477,WX9476);
  not NOT_3143(WX9480,WX10054);
  not NOT_3144(WX9484,WX10055);
  not NOT_3145(WX9488,WX10055);
  not NOT_3146(WX9490,WX9481);
  not NOT_3147(WX9491,WX9490);
  not NOT_3148(WX9494,WX10054);
  not NOT_3149(WX9498,WX10055);
  not NOT_3150(WX9502,WX10055);
  not NOT_3151(WX9504,WX9495);
  not NOT_3152(WX9505,WX9504);
  not NOT_3153(WX9508,WX10054);
  not NOT_3154(WX9512,WX10055);
  not NOT_3155(WX9516,WX10055);
  not NOT_3156(WX9518,WX9509);
  not NOT_3157(WX9519,WX9518);
  not NOT_3158(WX9522,WX10054);
  not NOT_3159(WX9526,WX10055);
  not NOT_3160(WX9530,WX10055);
  not NOT_3161(WX9532,WX9523);
  not NOT_3162(WX9533,WX9532);
  not NOT_3163(WX9534,WX9536);
  not NOT_3164(WX9599,WX10016);
  not NOT_3165(WX9600,WX10018);
  not NOT_3166(WX9601,WX10020);
  not NOT_3167(WX9602,WX10022);
  not NOT_3168(WX9603,WX10024);
  not NOT_3169(WX9604,WX10026);
  not NOT_3170(WX9605,WX10028);
  not NOT_3171(WX9606,WX10030);
  not NOT_3172(WX9607,WX10032);
  not NOT_3173(WX9608,WX10034);
  not NOT_3174(WX9609,WX10036);
  not NOT_3175(WX9610,WX10038);
  not NOT_3176(WX9611,WX10040);
  not NOT_3177(WX9612,WX10042);
  not NOT_3178(WX9613,WX10044);
  not NOT_3179(WX9614,WX10046);
  not NOT_3180(WX9615,WX9984);
  not NOT_3181(WX9616,WX9986);
  not NOT_3182(WX9617,WX9988);
  not NOT_3183(WX9618,WX9990);
  not NOT_3184(WX9619,WX9992);
  not NOT_3185(WX9620,WX9994);
  not NOT_3186(WX9621,WX9996);
  not NOT_3187(WX9622,WX9998);
  not NOT_3188(WX9623,WX10000);
  not NOT_3189(WX9624,WX10002);
  not NOT_3190(WX9625,WX10004);
  not NOT_3191(WX9626,WX10006);
  not NOT_3192(WX9627,WX10008);
  not NOT_3193(WX9628,WX10010);
  not NOT_3194(WX9629,WX10012);
  not NOT_3195(WX9630,WX10014);
  not NOT_3196(WX9631,WX9599);
  not NOT_3197(WX9632,WX9600);
  not NOT_3198(WX9633,WX9601);
  not NOT_3199(WX9634,WX9602);
  not NOT_3200(WX9635,WX9603);
  not NOT_3201(WX9636,WX9604);
  not NOT_3202(WX9637,WX9605);
  not NOT_3203(WX9638,WX9606);
  not NOT_3204(WX9639,WX9607);
  not NOT_3205(WX9640,WX9608);
  not NOT_3206(WX9641,WX9609);
  not NOT_3207(WX9642,WX9610);
  not NOT_3208(WX9643,WX9611);
  not NOT_3209(WX9644,WX9612);
  not NOT_3210(WX9645,WX9613);
  not NOT_3211(WX9646,WX9614);
  not NOT_3212(WX9647,WX9615);
  not NOT_3213(WX9648,WX9616);
  not NOT_3214(WX9649,WX9617);
  not NOT_3215(WX9650,WX9618);
  not NOT_3216(WX9651,WX9619);
  not NOT_3217(WX9652,WX9620);
  not NOT_3218(WX9653,WX9621);
  not NOT_3219(WX9654,WX9622);
  not NOT_3220(WX9655,WX9623);
  not NOT_3221(WX9656,WX9624);
  not NOT_3222(WX9657,WX9625);
  not NOT_3223(WX9658,WX9626);
  not NOT_3224(WX9659,WX9627);
  not NOT_3225(WX9660,WX9628);
  not NOT_3226(WX9661,WX9629);
  not NOT_3227(WX9662,WX9630);
  not NOT_3228(WX9663,WX9888);
  not NOT_3229(WX9664,WX9890);
  not NOT_3230(WX9665,WX9892);
  not NOT_3231(WX9666,WX9894);
  not NOT_3232(WX9667,WX9896);
  not NOT_3233(WX9668,WX9898);
  not NOT_3234(WX9669,WX9900);
  not NOT_3235(WX9670,WX9902);
  not NOT_3236(WX9671,WX9904);
  not NOT_3237(WX9672,WX9906);
  not NOT_3238(WX9673,WX9908);
  not NOT_3239(WX9674,WX9910);
  not NOT_3240(WX9675,WX9912);
  not NOT_3241(WX9676,WX9914);
  not NOT_3242(WX9677,WX9916);
  not NOT_3243(WX9678,WX9918);
  not NOT_3244(WX9679,WX9920);
  not NOT_3245(WX9680,WX9922);
  not NOT_3246(WX9681,WX9924);
  not NOT_3247(WX9682,WX9926);
  not NOT_3248(WX9683,WX9928);
  not NOT_3249(WX9684,WX9930);
  not NOT_3250(WX9685,WX9932);
  not NOT_3251(WX9686,WX9934);
  not NOT_3252(WX9687,WX9936);
  not NOT_3253(WX9688,WX9938);
  not NOT_3254(WX9689,WX9940);
  not NOT_3255(WX9690,WX9942);
  not NOT_3256(WX9691,WX9944);
  not NOT_3257(WX9692,WX9946);
  not NOT_3258(WX9693,WX9948);
  not NOT_3259(WX9694,WX9950);
  not NOT_3260(WX9983,WX9967);
  not NOT_3261(WX9984,WX9983);
  not NOT_3262(WX9985,WX9968);
  not NOT_3263(WX9986,WX9985);
  not NOT_3264(WX9987,WX9969);
  not NOT_3265(WX9988,WX9987);
  not NOT_3266(WX9989,WX9970);
  not NOT_3267(WX9990,WX9989);
  not NOT_3268(WX9991,WX9971);
  not NOT_3269(WX9992,WX9991);
  not NOT_3270(WX9993,WX9972);
  not NOT_3271(WX9994,WX9993);
  not NOT_3272(WX9995,WX9973);
  not NOT_3273(WX9996,WX9995);
  not NOT_3274(WX9997,WX9974);
  not NOT_3275(WX9998,WX9997);
  not NOT_3276(WX9999,WX9975);
  not NOT_3277(WX10000,WX9999);
  not NOT_3278(WX10001,WX9976);
  not NOT_3279(WX10002,WX10001);
  not NOT_3280(WX10003,WX9977);
  not NOT_3281(WX10004,WX10003);
  not NOT_3282(WX10005,WX9978);
  not NOT_3283(WX10006,WX10005);
  not NOT_3284(WX10007,WX9979);
  not NOT_3285(WX10008,WX10007);
  not NOT_3286(WX10009,WX9980);
  not NOT_3287(WX10010,WX10009);
  not NOT_3288(WX10011,WX9981);
  not NOT_3289(WX10012,WX10011);
  not NOT_3290(WX10013,WX9982);
  not NOT_3291(WX10014,WX10013);
  not NOT_3292(WX10015,WX9951);
  not NOT_3293(WX10016,WX10015);
  not NOT_3294(WX10017,WX9952);
  not NOT_3295(WX10018,WX10017);
  not NOT_3296(WX10019,WX9953);
  not NOT_3297(WX10020,WX10019);
  not NOT_3298(WX10021,WX9954);
  not NOT_3299(WX10022,WX10021);
  not NOT_3300(WX10023,WX9955);
  not NOT_3301(WX10024,WX10023);
  not NOT_3302(WX10025,WX9956);
  not NOT_3303(WX10026,WX10025);
  not NOT_3304(WX10027,WX9957);
  not NOT_3305(WX10028,WX10027);
  not NOT_3306(WX10029,WX9958);
  not NOT_3307(WX10030,WX10029);
  not NOT_3308(WX10031,WX9959);
  not NOT_3309(WX10032,WX10031);
  not NOT_3310(WX10033,WX9960);
  not NOT_3311(WX10034,WX10033);
  not NOT_3312(WX10035,WX9961);
  not NOT_3313(WX10036,WX10035);
  not NOT_3314(WX10037,WX9962);
  not NOT_3315(WX10038,WX10037);
  not NOT_3316(WX10039,WX9963);
  not NOT_3317(WX10040,WX10039);
  not NOT_3318(WX10041,WX9964);
  not NOT_3319(WX10042,WX10041);
  not NOT_3320(WX10043,WX9965);
  not NOT_3321(WX10044,WX10043);
  not NOT_3322(WX10045,WX9966);
  not NOT_3323(WX10046,WX10045);
  not NOT_3324(WX10047,TM0);
  not NOT_3325(WX10048,TM0);
  not NOT_3326(WX10049,TM0);
  not NOT_3327(WX10050,TM1);
  not NOT_3328(WX10051,TM1);
  not NOT_3329(WX10052,WX10051);
  not NOT_3330(WX10053,WX10049);
  not NOT_3331(WX10054,WX10050);
  not NOT_3332(WX10055,WX10048);
  not NOT_3333(WX10056,WX10047);
  not NOT_3334(WX10060,WX10056);
  not NOT_3335(WX10062,WX10061);
  not NOT_3336(WX10063,WX10062);
  not NOT_3337(WX10067,WX10056);
  not NOT_3338(WX10069,WX10068);
  not NOT_3339(WX10070,WX10069);
  not NOT_3340(WX10074,WX10056);
  not NOT_3341(WX10076,WX10075);
  not NOT_3342(WX10077,WX10076);
  not NOT_3343(WX10081,WX10056);
  not NOT_3344(WX10083,WX10082);
  not NOT_3345(WX10084,WX10083);
  not NOT_3346(WX10088,WX10056);
  not NOT_3347(WX10090,WX10089);
  not NOT_3348(WX10091,WX10090);
  not NOT_3349(WX10095,WX10056);
  not NOT_3350(WX10097,WX10096);
  not NOT_3351(WX10098,WX10097);
  not NOT_3352(WX10102,WX10056);
  not NOT_3353(WX10104,WX10103);
  not NOT_3354(WX10105,WX10104);
  not NOT_3355(WX10109,WX10056);
  not NOT_3356(WX10111,WX10110);
  not NOT_3357(WX10112,WX10111);
  not NOT_3358(WX10116,WX10056);
  not NOT_3359(WX10118,WX10117);
  not NOT_3360(WX10119,WX10118);
  not NOT_3361(WX10123,WX10056);
  not NOT_3362(WX10125,WX10124);
  not NOT_3363(WX10126,WX10125);
  not NOT_3364(WX10130,WX10056);
  not NOT_3365(WX10132,WX10131);
  not NOT_3366(WX10133,WX10132);
  not NOT_3367(WX10137,WX10056);
  not NOT_3368(WX10139,WX10138);
  not NOT_3369(WX10140,WX10139);
  not NOT_3370(WX10144,WX10056);
  not NOT_3371(WX10146,WX10145);
  not NOT_3372(WX10147,WX10146);
  not NOT_3373(WX10151,WX10056);
  not NOT_3374(WX10153,WX10152);
  not NOT_3375(WX10154,WX10153);
  not NOT_3376(WX10158,WX10056);
  not NOT_3377(WX10160,WX10159);
  not NOT_3378(WX10161,WX10160);
  not NOT_3379(WX10165,WX10056);
  not NOT_3380(WX10167,WX10166);
  not NOT_3381(WX10168,WX10167);
  not NOT_3382(WX10172,WX10056);
  not NOT_3383(WX10174,WX10173);
  not NOT_3384(WX10175,WX10174);
  not NOT_3385(WX10179,WX10056);
  not NOT_3386(WX10181,WX10180);
  not NOT_3387(WX10182,WX10181);
  not NOT_3388(WX10186,WX10056);
  not NOT_3389(WX10188,WX10187);
  not NOT_3390(WX10189,WX10188);
  not NOT_3391(WX10193,WX10056);
  not NOT_3392(WX10195,WX10194);
  not NOT_3393(WX10196,WX10195);
  not NOT_3394(WX10200,WX10056);
  not NOT_3395(WX10202,WX10201);
  not NOT_3396(WX10203,WX10202);
  not NOT_3397(WX10207,WX10056);
  not NOT_3398(WX10209,WX10208);
  not NOT_3399(WX10210,WX10209);
  not NOT_3400(WX10214,WX10056);
  not NOT_3401(WX10216,WX10215);
  not NOT_3402(WX10217,WX10216);
  not NOT_3403(WX10221,WX10056);
  not NOT_3404(WX10223,WX10222);
  not NOT_3405(WX10224,WX10223);
  not NOT_3406(WX10228,WX10056);
  not NOT_3407(WX10230,WX10229);
  not NOT_3408(WX10231,WX10230);
  not NOT_3409(WX10235,WX10056);
  not NOT_3410(WX10237,WX10236);
  not NOT_3411(WX10238,WX10237);
  not NOT_3412(WX10242,WX10056);
  not NOT_3413(WX10244,WX10243);
  not NOT_3414(WX10245,WX10244);
  not NOT_3415(WX10249,WX10056);
  not NOT_3416(WX10251,WX10250);
  not NOT_3417(WX10252,WX10251);
  not NOT_3418(WX10256,WX10056);
  not NOT_3419(WX10258,WX10257);
  not NOT_3420(WX10259,WX10258);
  not NOT_3421(WX10263,WX10056);
  not NOT_3422(WX10265,WX10264);
  not NOT_3423(WX10266,WX10265);
  not NOT_3424(WX10270,WX10056);
  not NOT_3425(WX10272,WX10271);
  not NOT_3426(WX10273,WX10272);
  not NOT_3427(WX10277,WX10056);
  not NOT_3428(WX10279,WX10278);
  not NOT_3429(WX10280,WX10279);
  not NOT_3430(WX10281,RESET);
  not NOT_3431(WX10314,WX10281);
  not NOT_3432(WX10381,WX11347);
  not NOT_3433(WX10385,WX11348);
  not NOT_3434(WX10389,WX11348);
  not NOT_3435(WX10391,WX10382);
  not NOT_3436(WX10392,WX10391);
  not NOT_3437(WX10395,WX11347);
  not NOT_3438(WX10399,WX11348);
  not NOT_3439(WX10403,WX11348);
  not NOT_3440(WX10405,WX10396);
  not NOT_3441(WX10406,WX10405);
  not NOT_3442(WX10409,WX11347);
  not NOT_3443(WX10413,WX11348);
  not NOT_3444(WX10417,WX11348);
  not NOT_3445(WX10419,WX10410);
  not NOT_3446(WX10420,WX10419);
  not NOT_3447(WX10423,WX11347);
  not NOT_3448(WX10427,WX11348);
  not NOT_3449(WX10431,WX11348);
  not NOT_3450(WX10433,WX10424);
  not NOT_3451(WX10434,WX10433);
  not NOT_3452(WX10437,WX11347);
  not NOT_3453(WX10441,WX11348);
  not NOT_3454(WX10445,WX11348);
  not NOT_3455(WX10447,WX10438);
  not NOT_3456(WX10448,WX10447);
  not NOT_3457(WX10451,WX11347);
  not NOT_3458(WX10455,WX11348);
  not NOT_3459(WX10459,WX11348);
  not NOT_3460(WX10461,WX10452);
  not NOT_3461(WX10462,WX10461);
  not NOT_3462(WX10465,WX11347);
  not NOT_3463(WX10469,WX11348);
  not NOT_3464(WX10473,WX11348);
  not NOT_3465(WX10475,WX10466);
  not NOT_3466(WX10476,WX10475);
  not NOT_3467(WX10479,WX11347);
  not NOT_3468(WX10483,WX11348);
  not NOT_3469(WX10487,WX11348);
  not NOT_3470(WX10489,WX10480);
  not NOT_3471(WX10490,WX10489);
  not NOT_3472(WX10493,WX11347);
  not NOT_3473(WX10497,WX11348);
  not NOT_3474(WX10501,WX11348);
  not NOT_3475(WX10503,WX10494);
  not NOT_3476(WX10504,WX10503);
  not NOT_3477(WX10507,WX11347);
  not NOT_3478(WX10511,WX11348);
  not NOT_3479(WX10515,WX11348);
  not NOT_3480(WX10517,WX10508);
  not NOT_3481(WX10518,WX10517);
  not NOT_3482(WX10521,WX11347);
  not NOT_3483(WX10525,WX11348);
  not NOT_3484(WX10529,WX11348);
  not NOT_3485(WX10531,WX10522);
  not NOT_3486(WX10532,WX10531);
  not NOT_3487(WX10535,WX11347);
  not NOT_3488(WX10539,WX11348);
  not NOT_3489(WX10543,WX11348);
  not NOT_3490(WX10545,WX10536);
  not NOT_3491(WX10546,WX10545);
  not NOT_3492(WX10549,WX11347);
  not NOT_3493(WX10553,WX11348);
  not NOT_3494(WX10557,WX11348);
  not NOT_3495(WX10559,WX10550);
  not NOT_3496(WX10560,WX10559);
  not NOT_3497(WX10563,WX11347);
  not NOT_3498(WX10567,WX11348);
  not NOT_3499(WX10571,WX11348);
  not NOT_3500(WX10573,WX10564);
  not NOT_3501(WX10574,WX10573);
  not NOT_3502(WX10577,WX11347);
  not NOT_3503(WX10581,WX11348);
  not NOT_3504(WX10585,WX11348);
  not NOT_3505(WX10587,WX10578);
  not NOT_3506(WX10588,WX10587);
  not NOT_3507(WX10591,WX11347);
  not NOT_3508(WX10595,WX11348);
  not NOT_3509(WX10599,WX11348);
  not NOT_3510(WX10601,WX10592);
  not NOT_3511(WX10602,WX10601);
  not NOT_3512(WX10605,WX11347);
  not NOT_3513(WX10609,WX11348);
  not NOT_3514(WX10613,WX11348);
  not NOT_3515(WX10615,WX10606);
  not NOT_3516(WX10616,WX10615);
  not NOT_3517(WX10619,WX11347);
  not NOT_3518(WX10623,WX11348);
  not NOT_3519(WX10627,WX11348);
  not NOT_3520(WX10629,WX10620);
  not NOT_3521(WX10630,WX10629);
  not NOT_3522(WX10633,WX11347);
  not NOT_3523(WX10637,WX11348);
  not NOT_3524(WX10641,WX11348);
  not NOT_3525(WX10643,WX10634);
  not NOT_3526(WX10644,WX10643);
  not NOT_3527(WX10647,WX11347);
  not NOT_3528(WX10651,WX11348);
  not NOT_3529(WX10655,WX11348);
  not NOT_3530(WX10657,WX10648);
  not NOT_3531(WX10658,WX10657);
  not NOT_3532(WX10661,WX11347);
  not NOT_3533(WX10665,WX11348);
  not NOT_3534(WX10669,WX11348);
  not NOT_3535(WX10671,WX10662);
  not NOT_3536(WX10672,WX10671);
  not NOT_3537(WX10675,WX11347);
  not NOT_3538(WX10679,WX11348);
  not NOT_3539(WX10683,WX11348);
  not NOT_3540(WX10685,WX10676);
  not NOT_3541(WX10686,WX10685);
  not NOT_3542(WX10689,WX11347);
  not NOT_3543(WX10693,WX11348);
  not NOT_3544(WX10697,WX11348);
  not NOT_3545(WX10699,WX10690);
  not NOT_3546(WX10700,WX10699);
  not NOT_3547(WX10703,WX11347);
  not NOT_3548(WX10707,WX11348);
  not NOT_3549(WX10711,WX11348);
  not NOT_3550(WX10713,WX10704);
  not NOT_3551(WX10714,WX10713);
  not NOT_3552(WX10717,WX11347);
  not NOT_3553(WX10721,WX11348);
  not NOT_3554(WX10725,WX11348);
  not NOT_3555(WX10727,WX10718);
  not NOT_3556(WX10728,WX10727);
  not NOT_3557(WX10731,WX11347);
  not NOT_3558(WX10735,WX11348);
  not NOT_3559(WX10739,WX11348);
  not NOT_3560(WX10741,WX10732);
  not NOT_3561(WX10742,WX10741);
  not NOT_3562(WX10745,WX11347);
  not NOT_3563(WX10749,WX11348);
  not NOT_3564(WX10753,WX11348);
  not NOT_3565(WX10755,WX10746);
  not NOT_3566(WX10756,WX10755);
  not NOT_3567(WX10759,WX11347);
  not NOT_3568(WX10763,WX11348);
  not NOT_3569(WX10767,WX11348);
  not NOT_3570(WX10769,WX10760);
  not NOT_3571(WX10770,WX10769);
  not NOT_3572(WX10773,WX11347);
  not NOT_3573(WX10777,WX11348);
  not NOT_3574(WX10781,WX11348);
  not NOT_3575(WX10783,WX10774);
  not NOT_3576(WX10784,WX10783);
  not NOT_3577(WX10787,WX11347);
  not NOT_3578(WX10791,WX11348);
  not NOT_3579(WX10795,WX11348);
  not NOT_3580(WX10797,WX10788);
  not NOT_3581(WX10798,WX10797);
  not NOT_3582(WX10801,WX11347);
  not NOT_3583(WX10805,WX11348);
  not NOT_3584(WX10809,WX11348);
  not NOT_3585(WX10811,WX10802);
  not NOT_3586(WX10812,WX10811);
  not NOT_3587(WX10815,WX11347);
  not NOT_3588(WX10819,WX11348);
  not NOT_3589(WX10823,WX11348);
  not NOT_3590(WX10825,WX10816);
  not NOT_3591(WX10826,WX10825);
  not NOT_3592(WX10827,WX10829);
  not NOT_3593(WX10892,WX11309);
  not NOT_3594(WX10893,WX11311);
  not NOT_3595(WX10894,WX11313);
  not NOT_3596(WX10895,WX11315);
  not NOT_3597(WX10896,WX11317);
  not NOT_3598(WX10897,WX11319);
  not NOT_3599(WX10898,WX11321);
  not NOT_3600(WX10899,WX11323);
  not NOT_3601(WX10900,WX11325);
  not NOT_3602(WX10901,WX11327);
  not NOT_3603(WX10902,WX11329);
  not NOT_3604(WX10903,WX11331);
  not NOT_3605(WX10904,WX11333);
  not NOT_3606(WX10905,WX11335);
  not NOT_3607(WX10906,WX11337);
  not NOT_3608(WX10907,WX11339);
  not NOT_3609(WX10908,WX11277);
  not NOT_3610(WX10909,WX11279);
  not NOT_3611(WX10910,WX11281);
  not NOT_3612(WX10911,WX11283);
  not NOT_3613(WX10912,WX11285);
  not NOT_3614(WX10913,WX11287);
  not NOT_3615(WX10914,WX11289);
  not NOT_3616(WX10915,WX11291);
  not NOT_3617(WX10916,WX11293);
  not NOT_3618(WX10917,WX11295);
  not NOT_3619(WX10918,WX11297);
  not NOT_3620(WX10919,WX11299);
  not NOT_3621(WX10920,WX11301);
  not NOT_3622(WX10921,WX11303);
  not NOT_3623(WX10922,WX11305);
  not NOT_3624(WX10923,WX11307);
  not NOT_3625(WX10924,WX10892);
  not NOT_3626(WX10925,WX10893);
  not NOT_3627(WX10926,WX10894);
  not NOT_3628(WX10927,WX10895);
  not NOT_3629(WX10928,WX10896);
  not NOT_3630(WX10929,WX10897);
  not NOT_3631(WX10930,WX10898);
  not NOT_3632(WX10931,WX10899);
  not NOT_3633(WX10932,WX10900);
  not NOT_3634(WX10933,WX10901);
  not NOT_3635(WX10934,WX10902);
  not NOT_3636(WX10935,WX10903);
  not NOT_3637(WX10936,WX10904);
  not NOT_3638(WX10937,WX10905);
  not NOT_3639(WX10938,WX10906);
  not NOT_3640(WX10939,WX10907);
  not NOT_3641(WX10940,WX10908);
  not NOT_3642(WX10941,WX10909);
  not NOT_3643(WX10942,WX10910);
  not NOT_3644(WX10943,WX10911);
  not NOT_3645(WX10944,WX10912);
  not NOT_3646(WX10945,WX10913);
  not NOT_3647(WX10946,WX10914);
  not NOT_3648(WX10947,WX10915);
  not NOT_3649(WX10948,WX10916);
  not NOT_3650(WX10949,WX10917);
  not NOT_3651(WX10950,WX10918);
  not NOT_3652(WX10951,WX10919);
  not NOT_3653(WX10952,WX10920);
  not NOT_3654(WX10953,WX10921);
  not NOT_3655(WX10954,WX10922);
  not NOT_3656(WX10955,WX10923);
  not NOT_3657(WX10956,WX11181);
  not NOT_3658(WX10957,WX11183);
  not NOT_3659(WX10958,WX11185);
  not NOT_3660(WX10959,WX11187);
  not NOT_3661(WX10960,WX11189);
  not NOT_3662(WX10961,WX11191);
  not NOT_3663(WX10962,WX11193);
  not NOT_3664(WX10963,WX11195);
  not NOT_3665(WX10964,WX11197);
  not NOT_3666(WX10965,WX11199);
  not NOT_3667(WX10966,WX11201);
  not NOT_3668(WX10967,WX11203);
  not NOT_3669(WX10968,WX11205);
  not NOT_3670(WX10969,WX11207);
  not NOT_3671(WX10970,WX11209);
  not NOT_3672(WX10971,WX11211);
  not NOT_3673(WX10972,WX11213);
  not NOT_3674(WX10973,WX11215);
  not NOT_3675(WX10974,WX11217);
  not NOT_3676(WX10975,WX11219);
  not NOT_3677(WX10976,WX11221);
  not NOT_3678(WX10977,WX11223);
  not NOT_3679(WX10978,WX11225);
  not NOT_3680(WX10979,WX11227);
  not NOT_3681(WX10980,WX11229);
  not NOT_3682(WX10981,WX11231);
  not NOT_3683(WX10982,WX11233);
  not NOT_3684(WX10983,WX11235);
  not NOT_3685(WX10984,WX11237);
  not NOT_3686(WX10985,WX11239);
  not NOT_3687(WX10986,WX11241);
  not NOT_3688(WX10987,WX11243);
  not NOT_3689(WX11276,WX11260);
  not NOT_3690(WX11277,WX11276);
  not NOT_3691(WX11278,WX11261);
  not NOT_3692(WX11279,WX11278);
  not NOT_3693(WX11280,WX11262);
  not NOT_3694(WX11281,WX11280);
  not NOT_3695(WX11282,WX11263);
  not NOT_3696(WX11283,WX11282);
  not NOT_3697(WX11284,WX11264);
  not NOT_3698(WX11285,WX11284);
  not NOT_3699(WX11286,WX11265);
  not NOT_3700(WX11287,WX11286);
  not NOT_3701(WX11288,WX11266);
  not NOT_3702(WX11289,WX11288);
  not NOT_3703(WX11290,WX11267);
  not NOT_3704(WX11291,WX11290);
  not NOT_3705(WX11292,WX11268);
  not NOT_3706(WX11293,WX11292);
  not NOT_3707(WX11294,WX11269);
  not NOT_3708(WX11295,WX11294);
  not NOT_3709(WX11296,WX11270);
  not NOT_3710(WX11297,WX11296);
  not NOT_3711(WX11298,WX11271);
  not NOT_3712(WX11299,WX11298);
  not NOT_3713(WX11300,WX11272);
  not NOT_3714(WX11301,WX11300);
  not NOT_3715(WX11302,WX11273);
  not NOT_3716(WX11303,WX11302);
  not NOT_3717(WX11304,WX11274);
  not NOT_3718(WX11305,WX11304);
  not NOT_3719(WX11306,WX11275);
  not NOT_3720(WX11307,WX11306);
  not NOT_3721(WX11308,WX11244);
  not NOT_3722(WX11309,WX11308);
  not NOT_3723(WX11310,WX11245);
  not NOT_3724(WX11311,WX11310);
  not NOT_3725(WX11312,WX11246);
  not NOT_3726(WX11313,WX11312);
  not NOT_3727(WX11314,WX11247);
  not NOT_3728(WX11315,WX11314);
  not NOT_3729(WX11316,WX11248);
  not NOT_3730(WX11317,WX11316);
  not NOT_3731(WX11318,WX11249);
  not NOT_3732(WX11319,WX11318);
  not NOT_3733(WX11320,WX11250);
  not NOT_3734(WX11321,WX11320);
  not NOT_3735(WX11322,WX11251);
  not NOT_3736(WX11323,WX11322);
  not NOT_3737(WX11324,WX11252);
  not NOT_3738(WX11325,WX11324);
  not NOT_3739(WX11326,WX11253);
  not NOT_3740(WX11327,WX11326);
  not NOT_3741(WX11328,WX11254);
  not NOT_3742(WX11329,WX11328);
  not NOT_3743(WX11330,WX11255);
  not NOT_3744(WX11331,WX11330);
  not NOT_3745(WX11332,WX11256);
  not NOT_3746(WX11333,WX11332);
  not NOT_3747(WX11334,WX11257);
  not NOT_3748(WX11335,WX11334);
  not NOT_3749(WX11336,WX11258);
  not NOT_3750(WX11337,WX11336);
  not NOT_3751(WX11338,WX11259);
  not NOT_3752(WX11339,WX11338);
  not NOT_3753(WX11340,TM0);
  not NOT_3754(WX11341,TM0);
  not NOT_3755(WX11342,TM0);
  not NOT_3756(WX11343,TM1);
  not NOT_3757(WX11344,TM1);
  not NOT_3758(WX11345,WX11344);
  not NOT_3759(WX11346,WX11342);
  not NOT_3760(WX11347,WX11343);
  not NOT_3761(WX11348,WX11341);
  not NOT_3762(WX11349,WX11340);
  not NOT_3763(WX11353,WX11349);
  not NOT_3764(WX11355,WX11354);
  not NOT_3765(WX11356,WX11355);
  not NOT_3766(WX11360,WX11349);
  not NOT_3767(WX11362,WX11361);
  not NOT_3768(WX11363,WX11362);
  not NOT_3769(WX11367,WX11349);
  not NOT_3770(WX11369,WX11368);
  not NOT_3771(WX11370,WX11369);
  not NOT_3772(WX11374,WX11349);
  not NOT_3773(WX11376,WX11375);
  not NOT_3774(WX11377,WX11376);
  not NOT_3775(WX11381,WX11349);
  not NOT_3776(WX11383,WX11382);
  not NOT_3777(WX11384,WX11383);
  not NOT_3778(WX11388,WX11349);
  not NOT_3779(WX11390,WX11389);
  not NOT_3780(WX11391,WX11390);
  not NOT_3781(WX11395,WX11349);
  not NOT_3782(WX11397,WX11396);
  not NOT_3783(WX11398,WX11397);
  not NOT_3784(WX11402,WX11349);
  not NOT_3785(WX11404,WX11403);
  not NOT_3786(WX11405,WX11404);
  not NOT_3787(WX11409,WX11349);
  not NOT_3788(WX11411,WX11410);
  not NOT_3789(WX11412,WX11411);
  not NOT_3790(WX11416,WX11349);
  not NOT_3791(WX11418,WX11417);
  not NOT_3792(WX11419,WX11418);
  not NOT_3793(WX11423,WX11349);
  not NOT_3794(WX11425,WX11424);
  not NOT_3795(WX11426,WX11425);
  not NOT_3796(WX11430,WX11349);
  not NOT_3797(WX11432,WX11431);
  not NOT_3798(WX11433,WX11432);
  not NOT_3799(WX11437,WX11349);
  not NOT_3800(WX11439,WX11438);
  not NOT_3801(WX11440,WX11439);
  not NOT_3802(WX11444,WX11349);
  not NOT_3803(WX11446,WX11445);
  not NOT_3804(WX11447,WX11446);
  not NOT_3805(WX11451,WX11349);
  not NOT_3806(WX11453,WX11452);
  not NOT_3807(WX11454,WX11453);
  not NOT_3808(WX11458,WX11349);
  not NOT_3809(WX11460,WX11459);
  not NOT_3810(WX11461,WX11460);
  not NOT_3811(WX11465,WX11349);
  not NOT_3812(WX11467,WX11466);
  not NOT_3813(WX11468,WX11467);
  not NOT_3814(WX11472,WX11349);
  not NOT_3815(WX11474,WX11473);
  not NOT_3816(WX11475,WX11474);
  not NOT_3817(WX11479,WX11349);
  not NOT_3818(WX11481,WX11480);
  not NOT_3819(WX11482,WX11481);
  not NOT_3820(WX11486,WX11349);
  not NOT_3821(WX11488,WX11487);
  not NOT_3822(WX11489,WX11488);
  not NOT_3823(WX11493,WX11349);
  not NOT_3824(WX11495,WX11494);
  not NOT_3825(WX11496,WX11495);
  not NOT_3826(WX11500,WX11349);
  not NOT_3827(WX11502,WX11501);
  not NOT_3828(WX11503,WX11502);
  not NOT_3829(WX11507,WX11349);
  not NOT_3830(WX11509,WX11508);
  not NOT_3831(WX11510,WX11509);
  not NOT_3832(WX11514,WX11349);
  not NOT_3833(WX11516,WX11515);
  not NOT_3834(WX11517,WX11516);
  not NOT_3835(WX11521,WX11349);
  not NOT_3836(WX11523,WX11522);
  not NOT_3837(WX11524,WX11523);
  not NOT_3838(WX11528,WX11349);
  not NOT_3839(WX11530,WX11529);
  not NOT_3840(WX11531,WX11530);
  not NOT_3841(WX11535,WX11349);
  not NOT_3842(WX11537,WX11536);
  not NOT_3843(WX11538,WX11537);
  not NOT_3844(WX11542,WX11349);
  not NOT_3845(WX11544,WX11543);
  not NOT_3846(WX11545,WX11544);
  not NOT_3847(WX11549,WX11349);
  not NOT_3848(WX11551,WX11550);
  not NOT_3849(WX11552,WX11551);
  not NOT_3850(WX11556,WX11349);
  not NOT_3851(WX11558,WX11557);
  not NOT_3852(WX11559,WX11558);
  not NOT_3853(WX11563,WX11349);
  not NOT_3854(WX11565,WX11564);
  not NOT_3855(WX11566,WX11565);
  not NOT_3856(WX11570,WX11349);
  not NOT_3857(WX11572,WX11571);
  not NOT_3858(WX11573,WX11572);
  not NOT_3859(WX11574,RESET);
  not NOT_3860(WX11607,WX11574);
  and AND2_0(WX35,WX46,WX1003);
  and AND2_1(WX36,WX42,WX37);
  and AND2_2(WX39,CRC_OUT_9_31,WX1004);
  and AND2_3(WX40,WX2305,WX41);
  and AND2_4(WX43,WX485,WX1004);
  and AND2_5(WX44,DATA_9_31,WX45);
  and AND2_6(WX49,WX60,WX1003);
  and AND2_7(WX50,WX56,WX51);
  and AND2_8(WX53,CRC_OUT_9_30,WX1004);
  and AND2_9(WX54,WX2312,WX55);
  and AND2_10(WX57,WX487,WX1004);
  and AND2_11(WX58,DATA_9_30,WX59);
  and AND2_12(WX63,WX74,WX1003);
  and AND2_13(WX64,WX70,WX65);
  and AND2_14(WX67,CRC_OUT_9_29,WX1004);
  and AND2_15(WX68,WX2319,WX69);
  and AND2_16(WX71,WX489,WX1004);
  and AND2_17(WX72,DATA_9_29,WX73);
  and AND2_18(WX77,WX88,WX1003);
  and AND2_19(WX78,WX84,WX79);
  and AND2_20(WX81,CRC_OUT_9_28,WX1004);
  and AND2_21(WX82,WX2326,WX83);
  and AND2_22(WX85,WX491,WX1004);
  and AND2_23(WX86,DATA_9_28,WX87);
  and AND2_24(WX91,WX102,WX1003);
  and AND2_25(WX92,WX98,WX93);
  and AND2_26(WX95,CRC_OUT_9_27,WX1004);
  and AND2_27(WX96,WX2333,WX97);
  and AND2_28(WX99,WX493,WX1004);
  and AND2_29(WX100,DATA_9_27,WX101);
  and AND2_30(WX105,WX116,WX1003);
  and AND2_31(WX106,WX112,WX107);
  and AND2_32(WX109,CRC_OUT_9_26,WX1004);
  and AND2_33(WX110,WX2340,WX111);
  and AND2_34(WX113,WX495,WX1004);
  and AND2_35(WX114,DATA_9_26,WX115);
  and AND2_36(WX119,WX130,WX1003);
  and AND2_37(WX120,WX126,WX121);
  and AND2_38(WX123,CRC_OUT_9_25,WX1004);
  and AND2_39(WX124,WX2347,WX125);
  and AND2_40(WX127,WX497,WX1004);
  and AND2_41(WX128,DATA_9_25,WX129);
  and AND2_42(WX133,WX144,WX1003);
  and AND2_43(WX134,WX140,WX135);
  and AND2_44(WX137,CRC_OUT_9_24,WX1004);
  and AND2_45(WX138,WX2354,WX139);
  and AND2_46(WX141,WX499,WX1004);
  and AND2_47(WX142,DATA_9_24,WX143);
  and AND2_48(WX147,WX158,WX1003);
  and AND2_49(WX148,WX154,WX149);
  and AND2_50(WX151,CRC_OUT_9_23,WX1004);
  and AND2_51(WX152,WX2361,WX153);
  and AND2_52(WX155,WX501,WX1004);
  and AND2_53(WX156,DATA_9_23,WX157);
  and AND2_54(WX161,WX172,WX1003);
  and AND2_55(WX162,WX168,WX163);
  and AND2_56(WX165,CRC_OUT_9_22,WX1004);
  and AND2_57(WX166,WX2368,WX167);
  and AND2_58(WX169,WX503,WX1004);
  and AND2_59(WX170,DATA_9_22,WX171);
  and AND2_60(WX175,WX186,WX1003);
  and AND2_61(WX176,WX182,WX177);
  and AND2_62(WX179,CRC_OUT_9_21,WX1004);
  and AND2_63(WX180,WX2375,WX181);
  and AND2_64(WX183,WX505,WX1004);
  and AND2_65(WX184,DATA_9_21,WX185);
  and AND2_66(WX189,WX200,WX1003);
  and AND2_67(WX190,WX196,WX191);
  and AND2_68(WX193,CRC_OUT_9_20,WX1004);
  and AND2_69(WX194,WX2382,WX195);
  and AND2_70(WX197,WX507,WX1004);
  and AND2_71(WX198,DATA_9_20,WX199);
  and AND2_72(WX203,WX214,WX1003);
  and AND2_73(WX204,WX210,WX205);
  and AND2_74(WX207,CRC_OUT_9_19,WX1004);
  and AND2_75(WX208,WX2389,WX209);
  and AND2_76(WX211,WX509,WX1004);
  and AND2_77(WX212,DATA_9_19,WX213);
  and AND2_78(WX217,WX228,WX1003);
  and AND2_79(WX218,WX224,WX219);
  and AND2_80(WX221,CRC_OUT_9_18,WX1004);
  and AND2_81(WX222,WX2396,WX223);
  and AND2_82(WX225,WX511,WX1004);
  and AND2_83(WX226,DATA_9_18,WX227);
  and AND2_84(WX231,WX242,WX1003);
  and AND2_85(WX232,WX238,WX233);
  and AND2_86(WX235,CRC_OUT_9_17,WX1004);
  and AND2_87(WX236,WX2403,WX237);
  and AND2_88(WX239,WX513,WX1004);
  and AND2_89(WX240,DATA_9_17,WX241);
  and AND2_90(WX245,WX256,WX1003);
  and AND2_91(WX246,WX252,WX247);
  and AND2_92(WX249,CRC_OUT_9_16,WX1004);
  and AND2_93(WX250,WX2410,WX251);
  and AND2_94(WX253,WX515,WX1004);
  and AND2_95(WX254,DATA_9_16,WX255);
  and AND2_96(WX259,WX270,WX1003);
  and AND2_97(WX260,WX266,WX261);
  and AND2_98(WX263,CRC_OUT_9_15,WX1004);
  and AND2_99(WX264,WX2417,WX265);
  and AND2_100(WX267,WX517,WX1004);
  and AND2_101(WX268,DATA_9_15,WX269);
  and AND2_102(WX273,WX284,WX1003);
  and AND2_103(WX274,WX280,WX275);
  and AND2_104(WX277,CRC_OUT_9_14,WX1004);
  and AND2_105(WX278,WX2424,WX279);
  and AND2_106(WX281,WX519,WX1004);
  and AND2_107(WX282,DATA_9_14,WX283);
  and AND2_108(WX287,WX298,WX1003);
  and AND2_109(WX288,WX294,WX289);
  and AND2_110(WX291,CRC_OUT_9_13,WX1004);
  and AND2_111(WX292,WX2431,WX293);
  and AND2_112(WX295,WX521,WX1004);
  and AND2_113(WX296,DATA_9_13,WX297);
  and AND2_114(WX301,WX312,WX1003);
  and AND2_115(WX302,WX308,WX303);
  and AND2_116(WX305,CRC_OUT_9_12,WX1004);
  and AND2_117(WX306,WX2438,WX307);
  and AND2_118(WX309,WX523,WX1004);
  and AND2_119(WX310,DATA_9_12,WX311);
  and AND2_120(WX315,WX326,WX1003);
  and AND2_121(WX316,WX322,WX317);
  and AND2_122(WX319,CRC_OUT_9_11,WX1004);
  and AND2_123(WX320,WX2445,WX321);
  and AND2_124(WX323,WX525,WX1004);
  and AND2_125(WX324,DATA_9_11,WX325);
  and AND2_126(WX329,WX340,WX1003);
  and AND2_127(WX330,WX336,WX331);
  and AND2_128(WX333,CRC_OUT_9_10,WX1004);
  and AND2_129(WX334,WX2452,WX335);
  and AND2_130(WX337,WX527,WX1004);
  and AND2_131(WX338,DATA_9_10,WX339);
  and AND2_132(WX343,WX354,WX1003);
  and AND2_133(WX344,WX350,WX345);
  and AND2_134(WX347,CRC_OUT_9_9,WX1004);
  and AND2_135(WX348,WX2459,WX349);
  and AND2_136(WX351,WX529,WX1004);
  and AND2_137(WX352,DATA_9_9,WX353);
  and AND2_138(WX357,WX368,WX1003);
  and AND2_139(WX358,WX364,WX359);
  and AND2_140(WX361,CRC_OUT_9_8,WX1004);
  and AND2_141(WX362,WX2466,WX363);
  and AND2_142(WX365,WX531,WX1004);
  and AND2_143(WX366,DATA_9_8,WX367);
  and AND2_144(WX371,WX382,WX1003);
  and AND2_145(WX372,WX378,WX373);
  and AND2_146(WX375,CRC_OUT_9_7,WX1004);
  and AND2_147(WX376,WX2473,WX377);
  and AND2_148(WX379,WX533,WX1004);
  and AND2_149(WX380,DATA_9_7,WX381);
  and AND2_150(WX385,WX396,WX1003);
  and AND2_151(WX386,WX392,WX387);
  and AND2_152(WX389,CRC_OUT_9_6,WX1004);
  and AND2_153(WX390,WX2480,WX391);
  and AND2_154(WX393,WX535,WX1004);
  and AND2_155(WX394,DATA_9_6,WX395);
  and AND2_156(WX399,WX410,WX1003);
  and AND2_157(WX400,WX406,WX401);
  and AND2_158(WX403,CRC_OUT_9_5,WX1004);
  and AND2_159(WX404,WX2487,WX405);
  and AND2_160(WX407,WX537,WX1004);
  and AND2_161(WX408,DATA_9_5,WX409);
  and AND2_162(WX413,WX424,WX1003);
  and AND2_163(WX414,WX420,WX415);
  and AND2_164(WX417,CRC_OUT_9_4,WX1004);
  and AND2_165(WX418,WX2494,WX419);
  and AND2_166(WX421,WX539,WX1004);
  and AND2_167(WX422,DATA_9_4,WX423);
  and AND2_168(WX427,WX438,WX1003);
  and AND2_169(WX428,WX434,WX429);
  and AND2_170(WX431,CRC_OUT_9_3,WX1004);
  and AND2_171(WX432,WX2501,WX433);
  and AND2_172(WX435,WX541,WX1004);
  and AND2_173(WX436,DATA_9_3,WX437);
  and AND2_174(WX441,WX452,WX1003);
  and AND2_175(WX442,WX448,WX443);
  and AND2_176(WX445,CRC_OUT_9_2,WX1004);
  and AND2_177(WX446,WX2508,WX447);
  and AND2_178(WX449,WX543,WX1004);
  and AND2_179(WX450,DATA_9_2,WX451);
  and AND2_180(WX455,WX466,WX1003);
  and AND2_181(WX456,WX462,WX457);
  and AND2_182(WX459,CRC_OUT_9_1,WX1004);
  and AND2_183(WX460,WX2515,WX461);
  and AND2_184(WX463,WX545,WX1004);
  and AND2_185(WX464,DATA_9_1,WX465);
  and AND2_186(WX469,WX480,WX1003);
  and AND2_187(WX470,WX476,WX471);
  and AND2_188(WX473,CRC_OUT_9_0,WX1004);
  and AND2_189(WX474,WX2522,WX475);
  and AND2_190(WX477,WX547,WX1004);
  and AND2_191(WX478,DATA_9_0,WX479);
  and AND2_192(WX484,WX487,RESET);
  and AND2_193(WX486,WX489,RESET);
  and AND2_194(WX488,WX491,RESET);
  and AND2_195(WX490,WX493,RESET);
  and AND2_196(WX492,WX495,RESET);
  and AND2_197(WX494,WX497,RESET);
  and AND2_198(WX496,WX499,RESET);
  and AND2_199(WX498,WX501,RESET);
  and AND2_200(WX500,WX503,RESET);
  and AND2_201(WX502,WX505,RESET);
  and AND2_202(WX504,WX507,RESET);
  and AND2_203(WX506,WX509,RESET);
  and AND2_204(WX508,WX511,RESET);
  and AND2_205(WX510,WX513,RESET);
  and AND2_206(WX512,WX515,RESET);
  and AND2_207(WX514,WX517,RESET);
  and AND2_208(WX516,WX519,RESET);
  and AND2_209(WX518,WX521,RESET);
  and AND2_210(WX520,WX523,RESET);
  and AND2_211(WX522,WX525,RESET);
  and AND2_212(WX524,WX527,RESET);
  and AND2_213(WX526,WX529,RESET);
  and AND2_214(WX528,WX531,RESET);
  and AND2_215(WX530,WX533,RESET);
  and AND2_216(WX532,WX535,RESET);
  and AND2_217(WX534,WX537,RESET);
  and AND2_218(WX536,WX539,RESET);
  and AND2_219(WX538,WX541,RESET);
  and AND2_220(WX540,WX543,RESET);
  and AND2_221(WX542,WX545,RESET);
  and AND2_222(WX544,WX547,RESET);
  and AND2_223(WX546,WX483,RESET);
  and AND2_224(WX644,WX48,RESET);
  and AND2_225(WX646,WX62,RESET);
  and AND2_226(WX648,WX76,RESET);
  and AND2_227(WX650,WX90,RESET);
  and AND2_228(WX652,WX104,RESET);
  and AND2_229(WX654,WX118,RESET);
  and AND2_230(WX656,WX132,RESET);
  and AND2_231(WX658,WX146,RESET);
  and AND2_232(WX660,WX160,RESET);
  and AND2_233(WX662,WX174,RESET);
  and AND2_234(WX664,WX188,RESET);
  and AND2_235(WX666,WX202,RESET);
  and AND2_236(WX668,WX216,RESET);
  and AND2_237(WX670,WX230,RESET);
  and AND2_238(WX672,WX244,RESET);
  and AND2_239(WX674,WX258,RESET);
  and AND2_240(WX676,WX272,RESET);
  and AND2_241(WX678,WX286,RESET);
  and AND2_242(WX680,WX300,RESET);
  and AND2_243(WX682,WX314,RESET);
  and AND2_244(WX684,WX328,RESET);
  and AND2_245(WX686,WX342,RESET);
  and AND2_246(WX688,WX356,RESET);
  and AND2_247(WX690,WX370,RESET);
  and AND2_248(WX692,WX384,RESET);
  and AND2_249(WX694,WX398,RESET);
  and AND2_250(WX696,WX412,RESET);
  and AND2_251(WX698,WX426,RESET);
  and AND2_252(WX700,WX440,RESET);
  and AND2_253(WX702,WX454,RESET);
  and AND2_254(WX704,WX468,RESET);
  and AND2_255(WX706,WX482,RESET);
  and AND2_256(WX708,WX645,RESET);
  and AND2_257(WX710,WX647,RESET);
  and AND2_258(WX712,WX649,RESET);
  and AND2_259(WX714,WX651,RESET);
  and AND2_260(WX716,WX653,RESET);
  and AND2_261(WX718,WX655,RESET);
  and AND2_262(WX720,WX657,RESET);
  and AND2_263(WX722,WX659,RESET);
  and AND2_264(WX724,WX661,RESET);
  and AND2_265(WX726,WX663,RESET);
  and AND2_266(WX728,WX665,RESET);
  and AND2_267(WX730,WX667,RESET);
  and AND2_268(WX732,WX669,RESET);
  and AND2_269(WX734,WX671,RESET);
  and AND2_270(WX736,WX673,RESET);
  and AND2_271(WX738,WX675,RESET);
  and AND2_272(WX740,WX677,RESET);
  and AND2_273(WX742,WX679,RESET);
  and AND2_274(WX744,WX681,RESET);
  and AND2_275(WX746,WX683,RESET);
  and AND2_276(WX748,WX685,RESET);
  and AND2_277(WX750,WX687,RESET);
  and AND2_278(WX752,WX689,RESET);
  and AND2_279(WX754,WX691,RESET);
  and AND2_280(WX756,WX693,RESET);
  and AND2_281(WX758,WX695,RESET);
  and AND2_282(WX760,WX697,RESET);
  and AND2_283(WX762,WX699,RESET);
  and AND2_284(WX764,WX701,RESET);
  and AND2_285(WX766,WX703,RESET);
  and AND2_286(WX768,WX705,RESET);
  and AND2_287(WX770,WX707,RESET);
  and AND2_288(WX772,WX709,RESET);
  and AND2_289(WX774,WX711,RESET);
  and AND2_290(WX776,WX713,RESET);
  and AND2_291(WX778,WX715,RESET);
  and AND2_292(WX780,WX717,RESET);
  and AND2_293(WX782,WX719,RESET);
  and AND2_294(WX784,WX721,RESET);
  and AND2_295(WX786,WX723,RESET);
  and AND2_296(WX788,WX725,RESET);
  and AND2_297(WX790,WX727,RESET);
  and AND2_298(WX792,WX729,RESET);
  and AND2_299(WX794,WX731,RESET);
  and AND2_300(WX796,WX733,RESET);
  and AND2_301(WX798,WX735,RESET);
  and AND2_302(WX800,WX737,RESET);
  and AND2_303(WX802,WX739,RESET);
  and AND2_304(WX804,WX741,RESET);
  and AND2_305(WX806,WX743,RESET);
  and AND2_306(WX808,WX745,RESET);
  and AND2_307(WX810,WX747,RESET);
  and AND2_308(WX812,WX749,RESET);
  and AND2_309(WX814,WX751,RESET);
  and AND2_310(WX816,WX753,RESET);
  and AND2_311(WX818,WX755,RESET);
  and AND2_312(WX820,WX757,RESET);
  and AND2_313(WX822,WX759,RESET);
  and AND2_314(WX824,WX761,RESET);
  and AND2_315(WX826,WX763,RESET);
  and AND2_316(WX828,WX765,RESET);
  and AND2_317(WX830,WX767,RESET);
  and AND2_318(WX832,WX769,RESET);
  and AND2_319(WX834,WX771,RESET);
  and AND2_320(WX836,WX773,RESET);
  and AND2_321(WX838,WX775,RESET);
  and AND2_322(WX840,WX777,RESET);
  and AND2_323(WX842,WX779,RESET);
  and AND2_324(WX844,WX781,RESET);
  and AND2_325(WX846,WX783,RESET);
  and AND2_326(WX848,WX785,RESET);
  and AND2_327(WX850,WX787,RESET);
  and AND2_328(WX852,WX789,RESET);
  and AND2_329(WX854,WX791,RESET);
  and AND2_330(WX856,WX793,RESET);
  and AND2_331(WX858,WX795,RESET);
  and AND2_332(WX860,WX797,RESET);
  and AND2_333(WX862,WX799,RESET);
  and AND2_334(WX864,WX801,RESET);
  and AND2_335(WX866,WX803,RESET);
  and AND2_336(WX868,WX805,RESET);
  and AND2_337(WX870,WX807,RESET);
  and AND2_338(WX872,WX809,RESET);
  and AND2_339(WX874,WX811,RESET);
  and AND2_340(WX876,WX813,RESET);
  and AND2_341(WX878,WX815,RESET);
  and AND2_342(WX880,WX817,RESET);
  and AND2_343(WX882,WX819,RESET);
  and AND2_344(WX884,WX821,RESET);
  and AND2_345(WX886,WX823,RESET);
  and AND2_346(WX888,WX825,RESET);
  and AND2_347(WX890,WX827,RESET);
  and AND2_348(WX892,WX829,RESET);
  and AND2_349(WX894,WX831,RESET);
  and AND2_350(WX896,WX833,RESET);
  and AND2_351(WX898,WX835,RESET);
  and AND2_352(WX1007,WX1006,WX1005);
  and AND2_353(WX1008,WX580,WX1009);
  and AND2_354(WX1014,WX1013,WX1005);
  and AND2_355(WX1015,WX581,WX1016);
  and AND2_356(WX1021,WX1020,WX1005);
  and AND2_357(WX1022,WX582,WX1023);
  and AND2_358(WX1028,WX1027,WX1005);
  and AND2_359(WX1029,WX583,WX1030);
  and AND2_360(WX1035,WX1034,WX1005);
  and AND2_361(WX1036,WX584,WX1037);
  and AND2_362(WX1042,WX1041,WX1005);
  and AND2_363(WX1043,WX585,WX1044);
  and AND2_364(WX1049,WX1048,WX1005);
  and AND2_365(WX1050,WX586,WX1051);
  and AND2_366(WX1056,WX1055,WX1005);
  and AND2_367(WX1057,WX587,WX1058);
  and AND2_368(WX1063,WX1062,WX1005);
  and AND2_369(WX1064,WX588,WX1065);
  and AND2_370(WX1070,WX1069,WX1005);
  and AND2_371(WX1071,WX589,WX1072);
  and AND2_372(WX1077,WX1076,WX1005);
  and AND2_373(WX1078,WX590,WX1079);
  and AND2_374(WX1084,WX1083,WX1005);
  and AND2_375(WX1085,WX591,WX1086);
  and AND2_376(WX1091,WX1090,WX1005);
  and AND2_377(WX1092,WX592,WX1093);
  and AND2_378(WX1098,WX1097,WX1005);
  and AND2_379(WX1099,WX593,WX1100);
  and AND2_380(WX1105,WX1104,WX1005);
  and AND2_381(WX1106,WX594,WX1107);
  and AND2_382(WX1112,WX1111,WX1005);
  and AND2_383(WX1113,WX595,WX1114);
  and AND2_384(WX1119,WX1118,WX1005);
  and AND2_385(WX1120,WX596,WX1121);
  and AND2_386(WX1126,WX1125,WX1005);
  and AND2_387(WX1127,WX597,WX1128);
  and AND2_388(WX1133,WX1132,WX1005);
  and AND2_389(WX1134,WX598,WX1135);
  and AND2_390(WX1140,WX1139,WX1005);
  and AND2_391(WX1141,WX599,WX1142);
  and AND2_392(WX1147,WX1146,WX1005);
  and AND2_393(WX1148,WX600,WX1149);
  and AND2_394(WX1154,WX1153,WX1005);
  and AND2_395(WX1155,WX601,WX1156);
  and AND2_396(WX1161,WX1160,WX1005);
  and AND2_397(WX1162,WX602,WX1163);
  and AND2_398(WX1168,WX1167,WX1005);
  and AND2_399(WX1169,WX603,WX1170);
  and AND2_400(WX1175,WX1174,WX1005);
  and AND2_401(WX1176,WX604,WX1177);
  and AND2_402(WX1182,WX1181,WX1005);
  and AND2_403(WX1183,WX605,WX1184);
  and AND2_404(WX1189,WX1188,WX1005);
  and AND2_405(WX1190,WX606,WX1191);
  and AND2_406(WX1196,WX1195,WX1005);
  and AND2_407(WX1197,WX607,WX1198);
  and AND2_408(WX1203,WX1202,WX1005);
  and AND2_409(WX1204,WX608,WX1205);
  and AND2_410(WX1210,WX1209,WX1005);
  and AND2_411(WX1211,WX609,WX1212);
  and AND2_412(WX1217,WX1216,WX1005);
  and AND2_413(WX1218,WX610,WX1219);
  and AND2_414(WX1224,WX1223,WX1005);
  and AND2_415(WX1225,WX611,WX1226);
  and AND2_416(WX1264,WX1234,WX1263);
  and AND2_417(WX1266,WX1262,WX1263);
  and AND2_418(WX1268,WX1261,WX1263);
  and AND2_419(WX1270,WX1260,WX1263);
  and AND2_420(WX1272,WX1233,WX1263);
  and AND2_421(WX1274,WX1259,WX1263);
  and AND2_422(WX1276,WX1258,WX1263);
  and AND2_423(WX1278,WX1257,WX1263);
  and AND2_424(WX1280,WX1256,WX1263);
  and AND2_425(WX1282,WX1255,WX1263);
  and AND2_426(WX1284,WX1254,WX1263);
  and AND2_427(WX1286,WX1232,WX1263);
  and AND2_428(WX1288,WX1253,WX1263);
  and AND2_429(WX1290,WX1252,WX1263);
  and AND2_430(WX1292,WX1251,WX1263);
  and AND2_431(WX1294,WX1250,WX1263);
  and AND2_432(WX1296,WX1231,WX1263);
  and AND2_433(WX1298,WX1249,WX1263);
  and AND2_434(WX1300,WX1248,WX1263);
  and AND2_435(WX1302,WX1247,WX1263);
  and AND2_436(WX1304,WX1246,WX1263);
  and AND2_437(WX1306,WX1245,WX1263);
  and AND2_438(WX1308,WX1244,WX1263);
  and AND2_439(WX1310,WX1243,WX1263);
  and AND2_440(WX1312,WX1242,WX1263);
  and AND2_441(WX1314,WX1241,WX1263);
  and AND2_442(WX1316,WX1240,WX1263);
  and AND2_443(WX1318,WX1239,WX1263);
  and AND2_444(WX1320,WX1238,WX1263);
  and AND2_445(WX1322,WX1237,WX1263);
  and AND2_446(WX1324,WX1236,WX1263);
  and AND2_447(WX1326,WX1235,WX1263);
  and AND2_448(WX1328,WX1339,WX2296);
  and AND2_449(WX1329,WX1335,WX1330);
  and AND2_450(WX1332,CRC_OUT_8_31,WX2297);
  and AND2_451(WX1333,WX3598,WX1334);
  and AND2_452(WX1336,WX1778,WX2297);
  and AND2_453(WX1337,WX2305,WX1338);
  and AND2_454(WX1342,WX1353,WX2296);
  and AND2_455(WX1343,WX1349,WX1344);
  and AND2_456(WX1346,CRC_OUT_8_30,WX2297);
  and AND2_457(WX1347,WX3605,WX1348);
  and AND2_458(WX1350,WX1780,WX2297);
  and AND2_459(WX1351,WX2312,WX1352);
  and AND2_460(WX1356,WX1367,WX2296);
  and AND2_461(WX1357,WX1363,WX1358);
  and AND2_462(WX1360,CRC_OUT_8_29,WX2297);
  and AND2_463(WX1361,WX3612,WX1362);
  and AND2_464(WX1364,WX1782,WX2297);
  and AND2_465(WX1365,WX2319,WX1366);
  and AND2_466(WX1370,WX1381,WX2296);
  and AND2_467(WX1371,WX1377,WX1372);
  and AND2_468(WX1374,CRC_OUT_8_28,WX2297);
  and AND2_469(WX1375,WX3619,WX1376);
  and AND2_470(WX1378,WX1784,WX2297);
  and AND2_471(WX1379,WX2326,WX1380);
  and AND2_472(WX1384,WX1395,WX2296);
  and AND2_473(WX1385,WX1391,WX1386);
  and AND2_474(WX1388,CRC_OUT_8_27,WX2297);
  and AND2_475(WX1389,WX3626,WX1390);
  and AND2_476(WX1392,WX1786,WX2297);
  and AND2_477(WX1393,WX2333,WX1394);
  and AND2_478(WX1398,WX1409,WX2296);
  and AND2_479(WX1399,WX1405,WX1400);
  and AND2_480(WX1402,CRC_OUT_8_26,WX2297);
  and AND2_481(WX1403,WX3633,WX1404);
  and AND2_482(WX1406,WX1788,WX2297);
  and AND2_483(WX1407,WX2340,WX1408);
  and AND2_484(WX1412,WX1423,WX2296);
  and AND2_485(WX1413,WX1419,WX1414);
  and AND2_486(WX1416,CRC_OUT_8_25,WX2297);
  and AND2_487(WX1417,WX3640,WX1418);
  and AND2_488(WX1420,WX1790,WX2297);
  and AND2_489(WX1421,WX2347,WX1422);
  and AND2_490(WX1426,WX1437,WX2296);
  and AND2_491(WX1427,WX1433,WX1428);
  and AND2_492(WX1430,CRC_OUT_8_24,WX2297);
  and AND2_493(WX1431,WX3647,WX1432);
  and AND2_494(WX1434,WX1792,WX2297);
  and AND2_495(WX1435,WX2354,WX1436);
  and AND2_496(WX1440,WX1451,WX2296);
  and AND2_497(WX1441,WX1447,WX1442);
  and AND2_498(WX1444,CRC_OUT_8_23,WX2297);
  and AND2_499(WX1445,WX3654,WX1446);
  and AND2_500(WX1448,WX1794,WX2297);
  and AND2_501(WX1449,WX2361,WX1450);
  and AND2_502(WX1454,WX1465,WX2296);
  and AND2_503(WX1455,WX1461,WX1456);
  and AND2_504(WX1458,CRC_OUT_8_22,WX2297);
  and AND2_505(WX1459,WX3661,WX1460);
  and AND2_506(WX1462,WX1796,WX2297);
  and AND2_507(WX1463,WX2368,WX1464);
  and AND2_508(WX1468,WX1479,WX2296);
  and AND2_509(WX1469,WX1475,WX1470);
  and AND2_510(WX1472,CRC_OUT_8_21,WX2297);
  and AND2_511(WX1473,WX3668,WX1474);
  and AND2_512(WX1476,WX1798,WX2297);
  and AND2_513(WX1477,WX2375,WX1478);
  and AND2_514(WX1482,WX1493,WX2296);
  and AND2_515(WX1483,WX1489,WX1484);
  and AND2_516(WX1486,CRC_OUT_8_20,WX2297);
  and AND2_517(WX1487,WX3675,WX1488);
  and AND2_518(WX1490,WX1800,WX2297);
  and AND2_519(WX1491,WX2382,WX1492);
  and AND2_520(WX1496,WX1507,WX2296);
  and AND2_521(WX1497,WX1503,WX1498);
  and AND2_522(WX1500,CRC_OUT_8_19,WX2297);
  and AND2_523(WX1501,WX3682,WX1502);
  and AND2_524(WX1504,WX1802,WX2297);
  and AND2_525(WX1505,WX2389,WX1506);
  and AND2_526(WX1510,WX1521,WX2296);
  and AND2_527(WX1511,WX1517,WX1512);
  and AND2_528(WX1514,CRC_OUT_8_18,WX2297);
  and AND2_529(WX1515,WX3689,WX1516);
  and AND2_530(WX1518,WX1804,WX2297);
  and AND2_531(WX1519,WX2396,WX1520);
  and AND2_532(WX1524,WX1535,WX2296);
  and AND2_533(WX1525,WX1531,WX1526);
  and AND2_534(WX1528,CRC_OUT_8_17,WX2297);
  and AND2_535(WX1529,WX3696,WX1530);
  and AND2_536(WX1532,WX1806,WX2297);
  and AND2_537(WX1533,WX2403,WX1534);
  and AND2_538(WX1538,WX1549,WX2296);
  and AND2_539(WX1539,WX1545,WX1540);
  and AND2_540(WX1542,CRC_OUT_8_16,WX2297);
  and AND2_541(WX1543,WX3703,WX1544);
  and AND2_542(WX1546,WX1808,WX2297);
  and AND2_543(WX1547,WX2410,WX1548);
  and AND2_544(WX1552,WX1563,WX2296);
  and AND2_545(WX1553,WX1559,WX1554);
  and AND2_546(WX1556,CRC_OUT_8_15,WX2297);
  and AND2_547(WX1557,WX3710,WX1558);
  and AND2_548(WX1560,WX1810,WX2297);
  and AND2_549(WX1561,WX2417,WX1562);
  and AND2_550(WX1566,WX1577,WX2296);
  and AND2_551(WX1567,WX1573,WX1568);
  and AND2_552(WX1570,CRC_OUT_8_14,WX2297);
  and AND2_553(WX1571,WX3717,WX1572);
  and AND2_554(WX1574,WX1812,WX2297);
  and AND2_555(WX1575,WX2424,WX1576);
  and AND2_556(WX1580,WX1591,WX2296);
  and AND2_557(WX1581,WX1587,WX1582);
  and AND2_558(WX1584,CRC_OUT_8_13,WX2297);
  and AND2_559(WX1585,WX3724,WX1586);
  and AND2_560(WX1588,WX1814,WX2297);
  and AND2_561(WX1589,WX2431,WX1590);
  and AND2_562(WX1594,WX1605,WX2296);
  and AND2_563(WX1595,WX1601,WX1596);
  and AND2_564(WX1598,CRC_OUT_8_12,WX2297);
  and AND2_565(WX1599,WX3731,WX1600);
  and AND2_566(WX1602,WX1816,WX2297);
  and AND2_567(WX1603,WX2438,WX1604);
  and AND2_568(WX1608,WX1619,WX2296);
  and AND2_569(WX1609,WX1615,WX1610);
  and AND2_570(WX1612,CRC_OUT_8_11,WX2297);
  and AND2_571(WX1613,WX3738,WX1614);
  and AND2_572(WX1616,WX1818,WX2297);
  and AND2_573(WX1617,WX2445,WX1618);
  and AND2_574(WX1622,WX1633,WX2296);
  and AND2_575(WX1623,WX1629,WX1624);
  and AND2_576(WX1626,CRC_OUT_8_10,WX2297);
  and AND2_577(WX1627,WX3745,WX1628);
  and AND2_578(WX1630,WX1820,WX2297);
  and AND2_579(WX1631,WX2452,WX1632);
  and AND2_580(WX1636,WX1647,WX2296);
  and AND2_581(WX1637,WX1643,WX1638);
  and AND2_582(WX1640,CRC_OUT_8_9,WX2297);
  and AND2_583(WX1641,WX3752,WX1642);
  and AND2_584(WX1644,WX1822,WX2297);
  and AND2_585(WX1645,WX2459,WX1646);
  and AND2_586(WX1650,WX1661,WX2296);
  and AND2_587(WX1651,WX1657,WX1652);
  and AND2_588(WX1654,CRC_OUT_8_8,WX2297);
  and AND2_589(WX1655,WX3759,WX1656);
  and AND2_590(WX1658,WX1824,WX2297);
  and AND2_591(WX1659,WX2466,WX1660);
  and AND2_592(WX1664,WX1675,WX2296);
  and AND2_593(WX1665,WX1671,WX1666);
  and AND2_594(WX1668,CRC_OUT_8_7,WX2297);
  and AND2_595(WX1669,WX3766,WX1670);
  and AND2_596(WX1672,WX1826,WX2297);
  and AND2_597(WX1673,WX2473,WX1674);
  and AND2_598(WX1678,WX1689,WX2296);
  and AND2_599(WX1679,WX1685,WX1680);
  and AND2_600(WX1682,CRC_OUT_8_6,WX2297);
  and AND2_601(WX1683,WX3773,WX1684);
  and AND2_602(WX1686,WX1828,WX2297);
  and AND2_603(WX1687,WX2480,WX1688);
  and AND2_604(WX1692,WX1703,WX2296);
  and AND2_605(WX1693,WX1699,WX1694);
  and AND2_606(WX1696,CRC_OUT_8_5,WX2297);
  and AND2_607(WX1697,WX3780,WX1698);
  and AND2_608(WX1700,WX1830,WX2297);
  and AND2_609(WX1701,WX2487,WX1702);
  and AND2_610(WX1706,WX1717,WX2296);
  and AND2_611(WX1707,WX1713,WX1708);
  and AND2_612(WX1710,CRC_OUT_8_4,WX2297);
  and AND2_613(WX1711,WX3787,WX1712);
  and AND2_614(WX1714,WX1832,WX2297);
  and AND2_615(WX1715,WX2494,WX1716);
  and AND2_616(WX1720,WX1731,WX2296);
  and AND2_617(WX1721,WX1727,WX1722);
  and AND2_618(WX1724,CRC_OUT_8_3,WX2297);
  and AND2_619(WX1725,WX3794,WX1726);
  and AND2_620(WX1728,WX1834,WX2297);
  and AND2_621(WX1729,WX2501,WX1730);
  and AND2_622(WX1734,WX1745,WX2296);
  and AND2_623(WX1735,WX1741,WX1736);
  and AND2_624(WX1738,CRC_OUT_8_2,WX2297);
  and AND2_625(WX1739,WX3801,WX1740);
  and AND2_626(WX1742,WX1836,WX2297);
  and AND2_627(WX1743,WX2508,WX1744);
  and AND2_628(WX1748,WX1759,WX2296);
  and AND2_629(WX1749,WX1755,WX1750);
  and AND2_630(WX1752,CRC_OUT_8_1,WX2297);
  and AND2_631(WX1753,WX3808,WX1754);
  and AND2_632(WX1756,WX1838,WX2297);
  and AND2_633(WX1757,WX2515,WX1758);
  and AND2_634(WX1762,WX1773,WX2296);
  and AND2_635(WX1763,WX1769,WX1764);
  and AND2_636(WX1766,CRC_OUT_8_0,WX2297);
  and AND2_637(WX1767,WX3815,WX1768);
  and AND2_638(WX1770,WX1840,WX2297);
  and AND2_639(WX1771,WX2522,WX1772);
  and AND2_640(WX1777,WX1780,RESET);
  and AND2_641(WX1779,WX1782,RESET);
  and AND2_642(WX1781,WX1784,RESET);
  and AND2_643(WX1783,WX1786,RESET);
  and AND2_644(WX1785,WX1788,RESET);
  and AND2_645(WX1787,WX1790,RESET);
  and AND2_646(WX1789,WX1792,RESET);
  and AND2_647(WX1791,WX1794,RESET);
  and AND2_648(WX1793,WX1796,RESET);
  and AND2_649(WX1795,WX1798,RESET);
  and AND2_650(WX1797,WX1800,RESET);
  and AND2_651(WX1799,WX1802,RESET);
  and AND2_652(WX1801,WX1804,RESET);
  and AND2_653(WX1803,WX1806,RESET);
  and AND2_654(WX1805,WX1808,RESET);
  and AND2_655(WX1807,WX1810,RESET);
  and AND2_656(WX1809,WX1812,RESET);
  and AND2_657(WX1811,WX1814,RESET);
  and AND2_658(WX1813,WX1816,RESET);
  and AND2_659(WX1815,WX1818,RESET);
  and AND2_660(WX1817,WX1820,RESET);
  and AND2_661(WX1819,WX1822,RESET);
  and AND2_662(WX1821,WX1824,RESET);
  and AND2_663(WX1823,WX1826,RESET);
  and AND2_664(WX1825,WX1828,RESET);
  and AND2_665(WX1827,WX1830,RESET);
  and AND2_666(WX1829,WX1832,RESET);
  and AND2_667(WX1831,WX1834,RESET);
  and AND2_668(WX1833,WX1836,RESET);
  and AND2_669(WX1835,WX1838,RESET);
  and AND2_670(WX1837,WX1840,RESET);
  and AND2_671(WX1839,WX1776,RESET);
  and AND2_672(WX1937,WX1341,RESET);
  and AND2_673(WX1939,WX1355,RESET);
  and AND2_674(WX1941,WX1369,RESET);
  and AND2_675(WX1943,WX1383,RESET);
  and AND2_676(WX1945,WX1397,RESET);
  and AND2_677(WX1947,WX1411,RESET);
  and AND2_678(WX1949,WX1425,RESET);
  and AND2_679(WX1951,WX1439,RESET);
  and AND2_680(WX1953,WX1453,RESET);
  and AND2_681(WX1955,WX1467,RESET);
  and AND2_682(WX1957,WX1481,RESET);
  and AND2_683(WX1959,WX1495,RESET);
  and AND2_684(WX1961,WX1509,RESET);
  and AND2_685(WX1963,WX1523,RESET);
  and AND2_686(WX1965,WX1537,RESET);
  and AND2_687(WX1967,WX1551,RESET);
  and AND2_688(WX1969,WX1565,RESET);
  and AND2_689(WX1971,WX1579,RESET);
  and AND2_690(WX1973,WX1593,RESET);
  and AND2_691(WX1975,WX1607,RESET);
  and AND2_692(WX1977,WX1621,RESET);
  and AND2_693(WX1979,WX1635,RESET);
  and AND2_694(WX1981,WX1649,RESET);
  and AND2_695(WX1983,WX1663,RESET);
  and AND2_696(WX1985,WX1677,RESET);
  and AND2_697(WX1987,WX1691,RESET);
  and AND2_698(WX1989,WX1705,RESET);
  and AND2_699(WX1991,WX1719,RESET);
  and AND2_700(WX1993,WX1733,RESET);
  and AND2_701(WX1995,WX1747,RESET);
  and AND2_702(WX1997,WX1761,RESET);
  and AND2_703(WX1999,WX1775,RESET);
  and AND2_704(WX2001,WX1938,RESET);
  and AND2_705(WX2003,WX1940,RESET);
  and AND2_706(WX2005,WX1942,RESET);
  and AND2_707(WX2007,WX1944,RESET);
  and AND2_708(WX2009,WX1946,RESET);
  and AND2_709(WX2011,WX1948,RESET);
  and AND2_710(WX2013,WX1950,RESET);
  and AND2_711(WX2015,WX1952,RESET);
  and AND2_712(WX2017,WX1954,RESET);
  and AND2_713(WX2019,WX1956,RESET);
  and AND2_714(WX2021,WX1958,RESET);
  and AND2_715(WX2023,WX1960,RESET);
  and AND2_716(WX2025,WX1962,RESET);
  and AND2_717(WX2027,WX1964,RESET);
  and AND2_718(WX2029,WX1966,RESET);
  and AND2_719(WX2031,WX1968,RESET);
  and AND2_720(WX2033,WX1970,RESET);
  and AND2_721(WX2035,WX1972,RESET);
  and AND2_722(WX2037,WX1974,RESET);
  and AND2_723(WX2039,WX1976,RESET);
  and AND2_724(WX2041,WX1978,RESET);
  and AND2_725(WX2043,WX1980,RESET);
  and AND2_726(WX2045,WX1982,RESET);
  and AND2_727(WX2047,WX1984,RESET);
  and AND2_728(WX2049,WX1986,RESET);
  and AND2_729(WX2051,WX1988,RESET);
  and AND2_730(WX2053,WX1990,RESET);
  and AND2_731(WX2055,WX1992,RESET);
  and AND2_732(WX2057,WX1994,RESET);
  and AND2_733(WX2059,WX1996,RESET);
  and AND2_734(WX2061,WX1998,RESET);
  and AND2_735(WX2063,WX2000,RESET);
  and AND2_736(WX2065,WX2002,RESET);
  and AND2_737(WX2067,WX2004,RESET);
  and AND2_738(WX2069,WX2006,RESET);
  and AND2_739(WX2071,WX2008,RESET);
  and AND2_740(WX2073,WX2010,RESET);
  and AND2_741(WX2075,WX2012,RESET);
  and AND2_742(WX2077,WX2014,RESET);
  and AND2_743(WX2079,WX2016,RESET);
  and AND2_744(WX2081,WX2018,RESET);
  and AND2_745(WX2083,WX2020,RESET);
  and AND2_746(WX2085,WX2022,RESET);
  and AND2_747(WX2087,WX2024,RESET);
  and AND2_748(WX2089,WX2026,RESET);
  and AND2_749(WX2091,WX2028,RESET);
  and AND2_750(WX2093,WX2030,RESET);
  and AND2_751(WX2095,WX2032,RESET);
  and AND2_752(WX2097,WX2034,RESET);
  and AND2_753(WX2099,WX2036,RESET);
  and AND2_754(WX2101,WX2038,RESET);
  and AND2_755(WX2103,WX2040,RESET);
  and AND2_756(WX2105,WX2042,RESET);
  and AND2_757(WX2107,WX2044,RESET);
  and AND2_758(WX2109,WX2046,RESET);
  and AND2_759(WX2111,WX2048,RESET);
  and AND2_760(WX2113,WX2050,RESET);
  and AND2_761(WX2115,WX2052,RESET);
  and AND2_762(WX2117,WX2054,RESET);
  and AND2_763(WX2119,WX2056,RESET);
  and AND2_764(WX2121,WX2058,RESET);
  and AND2_765(WX2123,WX2060,RESET);
  and AND2_766(WX2125,WX2062,RESET);
  and AND2_767(WX2127,WX2064,RESET);
  and AND2_768(WX2129,WX2066,RESET);
  and AND2_769(WX2131,WX2068,RESET);
  and AND2_770(WX2133,WX2070,RESET);
  and AND2_771(WX2135,WX2072,RESET);
  and AND2_772(WX2137,WX2074,RESET);
  and AND2_773(WX2139,WX2076,RESET);
  and AND2_774(WX2141,WX2078,RESET);
  and AND2_775(WX2143,WX2080,RESET);
  and AND2_776(WX2145,WX2082,RESET);
  and AND2_777(WX2147,WX2084,RESET);
  and AND2_778(WX2149,WX2086,RESET);
  and AND2_779(WX2151,WX2088,RESET);
  and AND2_780(WX2153,WX2090,RESET);
  and AND2_781(WX2155,WX2092,RESET);
  and AND2_782(WX2157,WX2094,RESET);
  and AND2_783(WX2159,WX2096,RESET);
  and AND2_784(WX2161,WX2098,RESET);
  and AND2_785(WX2163,WX2100,RESET);
  and AND2_786(WX2165,WX2102,RESET);
  and AND2_787(WX2167,WX2104,RESET);
  and AND2_788(WX2169,WX2106,RESET);
  and AND2_789(WX2171,WX2108,RESET);
  and AND2_790(WX2173,WX2110,RESET);
  and AND2_791(WX2175,WX2112,RESET);
  and AND2_792(WX2177,WX2114,RESET);
  and AND2_793(WX2179,WX2116,RESET);
  and AND2_794(WX2181,WX2118,RESET);
  and AND2_795(WX2183,WX2120,RESET);
  and AND2_796(WX2185,WX2122,RESET);
  and AND2_797(WX2187,WX2124,RESET);
  and AND2_798(WX2189,WX2126,RESET);
  and AND2_799(WX2191,WX2128,RESET);
  and AND2_800(WX2300,WX2299,WX2298);
  and AND2_801(WX2301,WX1873,WX2302);
  and AND2_802(WX2307,WX2306,WX2298);
  and AND2_803(WX2308,WX1874,WX2309);
  and AND2_804(WX2314,WX2313,WX2298);
  and AND2_805(WX2315,WX1875,WX2316);
  and AND2_806(WX2321,WX2320,WX2298);
  and AND2_807(WX2322,WX1876,WX2323);
  and AND2_808(WX2328,WX2327,WX2298);
  and AND2_809(WX2329,WX1877,WX2330);
  and AND2_810(WX2335,WX2334,WX2298);
  and AND2_811(WX2336,WX1878,WX2337);
  and AND2_812(WX2342,WX2341,WX2298);
  and AND2_813(WX2343,WX1879,WX2344);
  and AND2_814(WX2349,WX2348,WX2298);
  and AND2_815(WX2350,WX1880,WX2351);
  and AND2_816(WX2356,WX2355,WX2298);
  and AND2_817(WX2357,WX1881,WX2358);
  and AND2_818(WX2363,WX2362,WX2298);
  and AND2_819(WX2364,WX1882,WX2365);
  and AND2_820(WX2370,WX2369,WX2298);
  and AND2_821(WX2371,WX1883,WX2372);
  and AND2_822(WX2377,WX2376,WX2298);
  and AND2_823(WX2378,WX1884,WX2379);
  and AND2_824(WX2384,WX2383,WX2298);
  and AND2_825(WX2385,WX1885,WX2386);
  and AND2_826(WX2391,WX2390,WX2298);
  and AND2_827(WX2392,WX1886,WX2393);
  and AND2_828(WX2398,WX2397,WX2298);
  and AND2_829(WX2399,WX1887,WX2400);
  and AND2_830(WX2405,WX2404,WX2298);
  and AND2_831(WX2406,WX1888,WX2407);
  and AND2_832(WX2412,WX2411,WX2298);
  and AND2_833(WX2413,WX1889,WX2414);
  and AND2_834(WX2419,WX2418,WX2298);
  and AND2_835(WX2420,WX1890,WX2421);
  and AND2_836(WX2426,WX2425,WX2298);
  and AND2_837(WX2427,WX1891,WX2428);
  and AND2_838(WX2433,WX2432,WX2298);
  and AND2_839(WX2434,WX1892,WX2435);
  and AND2_840(WX2440,WX2439,WX2298);
  and AND2_841(WX2441,WX1893,WX2442);
  and AND2_842(WX2447,WX2446,WX2298);
  and AND2_843(WX2448,WX1894,WX2449);
  and AND2_844(WX2454,WX2453,WX2298);
  and AND2_845(WX2455,WX1895,WX2456);
  and AND2_846(WX2461,WX2460,WX2298);
  and AND2_847(WX2462,WX1896,WX2463);
  and AND2_848(WX2468,WX2467,WX2298);
  and AND2_849(WX2469,WX1897,WX2470);
  and AND2_850(WX2475,WX2474,WX2298);
  and AND2_851(WX2476,WX1898,WX2477);
  and AND2_852(WX2482,WX2481,WX2298);
  and AND2_853(WX2483,WX1899,WX2484);
  and AND2_854(WX2489,WX2488,WX2298);
  and AND2_855(WX2490,WX1900,WX2491);
  and AND2_856(WX2496,WX2495,WX2298);
  and AND2_857(WX2497,WX1901,WX2498);
  and AND2_858(WX2503,WX2502,WX2298);
  and AND2_859(WX2504,WX1902,WX2505);
  and AND2_860(WX2510,WX2509,WX2298);
  and AND2_861(WX2511,WX1903,WX2512);
  and AND2_862(WX2517,WX2516,WX2298);
  and AND2_863(WX2518,WX1904,WX2519);
  and AND2_864(WX2557,WX2527,WX2556);
  and AND2_865(WX2559,WX2555,WX2556);
  and AND2_866(WX2561,WX2554,WX2556);
  and AND2_867(WX2563,WX2553,WX2556);
  and AND2_868(WX2565,WX2526,WX2556);
  and AND2_869(WX2567,WX2552,WX2556);
  and AND2_870(WX2569,WX2551,WX2556);
  and AND2_871(WX2571,WX2550,WX2556);
  and AND2_872(WX2573,WX2549,WX2556);
  and AND2_873(WX2575,WX2548,WX2556);
  and AND2_874(WX2577,WX2547,WX2556);
  and AND2_875(WX2579,WX2525,WX2556);
  and AND2_876(WX2581,WX2546,WX2556);
  and AND2_877(WX2583,WX2545,WX2556);
  and AND2_878(WX2585,WX2544,WX2556);
  and AND2_879(WX2587,WX2543,WX2556);
  and AND2_880(WX2589,WX2524,WX2556);
  and AND2_881(WX2591,WX2542,WX2556);
  and AND2_882(WX2593,WX2541,WX2556);
  and AND2_883(WX2595,WX2540,WX2556);
  and AND2_884(WX2597,WX2539,WX2556);
  and AND2_885(WX2599,WX2538,WX2556);
  and AND2_886(WX2601,WX2537,WX2556);
  and AND2_887(WX2603,WX2536,WX2556);
  and AND2_888(WX2605,WX2535,WX2556);
  and AND2_889(WX2607,WX2534,WX2556);
  and AND2_890(WX2609,WX2533,WX2556);
  and AND2_891(WX2611,WX2532,WX2556);
  and AND2_892(WX2613,WX2531,WX2556);
  and AND2_893(WX2615,WX2530,WX2556);
  and AND2_894(WX2617,WX2529,WX2556);
  and AND2_895(WX2619,WX2528,WX2556);
  and AND2_896(WX2621,WX2632,WX3589);
  and AND2_897(WX2622,WX2628,WX2623);
  and AND2_898(WX2625,CRC_OUT_7_31,WX3590);
  and AND2_899(WX2626,WX4891,WX2627);
  and AND2_900(WX2629,WX3071,WX3590);
  and AND2_901(WX2630,WX3598,WX2631);
  and AND2_902(WX2635,WX2646,WX3589);
  and AND2_903(WX2636,WX2642,WX2637);
  and AND2_904(WX2639,CRC_OUT_7_30,WX3590);
  and AND2_905(WX2640,WX4898,WX2641);
  and AND2_906(WX2643,WX3073,WX3590);
  and AND2_907(WX2644,WX3605,WX2645);
  and AND2_908(WX2649,WX2660,WX3589);
  and AND2_909(WX2650,WX2656,WX2651);
  and AND2_910(WX2653,CRC_OUT_7_29,WX3590);
  and AND2_911(WX2654,WX4905,WX2655);
  and AND2_912(WX2657,WX3075,WX3590);
  and AND2_913(WX2658,WX3612,WX2659);
  and AND2_914(WX2663,WX2674,WX3589);
  and AND2_915(WX2664,WX2670,WX2665);
  and AND2_916(WX2667,CRC_OUT_7_28,WX3590);
  and AND2_917(WX2668,WX4912,WX2669);
  and AND2_918(WX2671,WX3077,WX3590);
  and AND2_919(WX2672,WX3619,WX2673);
  and AND2_920(WX2677,WX2688,WX3589);
  and AND2_921(WX2678,WX2684,WX2679);
  and AND2_922(WX2681,CRC_OUT_7_27,WX3590);
  and AND2_923(WX2682,WX4919,WX2683);
  and AND2_924(WX2685,WX3079,WX3590);
  and AND2_925(WX2686,WX3626,WX2687);
  and AND2_926(WX2691,WX2702,WX3589);
  and AND2_927(WX2692,WX2698,WX2693);
  and AND2_928(WX2695,CRC_OUT_7_26,WX3590);
  and AND2_929(WX2696,WX4926,WX2697);
  and AND2_930(WX2699,WX3081,WX3590);
  and AND2_931(WX2700,WX3633,WX2701);
  and AND2_932(WX2705,WX2716,WX3589);
  and AND2_933(WX2706,WX2712,WX2707);
  and AND2_934(WX2709,CRC_OUT_7_25,WX3590);
  and AND2_935(WX2710,WX4933,WX2711);
  and AND2_936(WX2713,WX3083,WX3590);
  and AND2_937(WX2714,WX3640,WX2715);
  and AND2_938(WX2719,WX2730,WX3589);
  and AND2_939(WX2720,WX2726,WX2721);
  and AND2_940(WX2723,CRC_OUT_7_24,WX3590);
  and AND2_941(WX2724,WX4940,WX2725);
  and AND2_942(WX2727,WX3085,WX3590);
  and AND2_943(WX2728,WX3647,WX2729);
  and AND2_944(WX2733,WX2744,WX3589);
  and AND2_945(WX2734,WX2740,WX2735);
  and AND2_946(WX2737,CRC_OUT_7_23,WX3590);
  and AND2_947(WX2738,WX4947,WX2739);
  and AND2_948(WX2741,WX3087,WX3590);
  and AND2_949(WX2742,WX3654,WX2743);
  and AND2_950(WX2747,WX2758,WX3589);
  and AND2_951(WX2748,WX2754,WX2749);
  and AND2_952(WX2751,CRC_OUT_7_22,WX3590);
  and AND2_953(WX2752,WX4954,WX2753);
  and AND2_954(WX2755,WX3089,WX3590);
  and AND2_955(WX2756,WX3661,WX2757);
  and AND2_956(WX2761,WX2772,WX3589);
  and AND2_957(WX2762,WX2768,WX2763);
  and AND2_958(WX2765,CRC_OUT_7_21,WX3590);
  and AND2_959(WX2766,WX4961,WX2767);
  and AND2_960(WX2769,WX3091,WX3590);
  and AND2_961(WX2770,WX3668,WX2771);
  and AND2_962(WX2775,WX2786,WX3589);
  and AND2_963(WX2776,WX2782,WX2777);
  and AND2_964(WX2779,CRC_OUT_7_20,WX3590);
  and AND2_965(WX2780,WX4968,WX2781);
  and AND2_966(WX2783,WX3093,WX3590);
  and AND2_967(WX2784,WX3675,WX2785);
  and AND2_968(WX2789,WX2800,WX3589);
  and AND2_969(WX2790,WX2796,WX2791);
  and AND2_970(WX2793,CRC_OUT_7_19,WX3590);
  and AND2_971(WX2794,WX4975,WX2795);
  and AND2_972(WX2797,WX3095,WX3590);
  and AND2_973(WX2798,WX3682,WX2799);
  and AND2_974(WX2803,WX2814,WX3589);
  and AND2_975(WX2804,WX2810,WX2805);
  and AND2_976(WX2807,CRC_OUT_7_18,WX3590);
  and AND2_977(WX2808,WX4982,WX2809);
  and AND2_978(WX2811,WX3097,WX3590);
  and AND2_979(WX2812,WX3689,WX2813);
  and AND2_980(WX2817,WX2828,WX3589);
  and AND2_981(WX2818,WX2824,WX2819);
  and AND2_982(WX2821,CRC_OUT_7_17,WX3590);
  and AND2_983(WX2822,WX4989,WX2823);
  and AND2_984(WX2825,WX3099,WX3590);
  and AND2_985(WX2826,WX3696,WX2827);
  and AND2_986(WX2831,WX2842,WX3589);
  and AND2_987(WX2832,WX2838,WX2833);
  and AND2_988(WX2835,CRC_OUT_7_16,WX3590);
  and AND2_989(WX2836,WX4996,WX2837);
  and AND2_990(WX2839,WX3101,WX3590);
  and AND2_991(WX2840,WX3703,WX2841);
  and AND2_992(WX2845,WX2856,WX3589);
  and AND2_993(WX2846,WX2852,WX2847);
  and AND2_994(WX2849,CRC_OUT_7_15,WX3590);
  and AND2_995(WX2850,WX5003,WX2851);
  and AND2_996(WX2853,WX3103,WX3590);
  and AND2_997(WX2854,WX3710,WX2855);
  and AND2_998(WX2859,WX2870,WX3589);
  and AND2_999(WX2860,WX2866,WX2861);
  and AND2_1000(WX2863,CRC_OUT_7_14,WX3590);
  and AND2_1001(WX2864,WX5010,WX2865);
  and AND2_1002(WX2867,WX3105,WX3590);
  and AND2_1003(WX2868,WX3717,WX2869);
  and AND2_1004(WX2873,WX2884,WX3589);
  and AND2_1005(WX2874,WX2880,WX2875);
  and AND2_1006(WX2877,CRC_OUT_7_13,WX3590);
  and AND2_1007(WX2878,WX5017,WX2879);
  and AND2_1008(WX2881,WX3107,WX3590);
  and AND2_1009(WX2882,WX3724,WX2883);
  and AND2_1010(WX2887,WX2898,WX3589);
  and AND2_1011(WX2888,WX2894,WX2889);
  and AND2_1012(WX2891,CRC_OUT_7_12,WX3590);
  and AND2_1013(WX2892,WX5024,WX2893);
  and AND2_1014(WX2895,WX3109,WX3590);
  and AND2_1015(WX2896,WX3731,WX2897);
  and AND2_1016(WX2901,WX2912,WX3589);
  and AND2_1017(WX2902,WX2908,WX2903);
  and AND2_1018(WX2905,CRC_OUT_7_11,WX3590);
  and AND2_1019(WX2906,WX5031,WX2907);
  and AND2_1020(WX2909,WX3111,WX3590);
  and AND2_1021(WX2910,WX3738,WX2911);
  and AND2_1022(WX2915,WX2926,WX3589);
  and AND2_1023(WX2916,WX2922,WX2917);
  and AND2_1024(WX2919,CRC_OUT_7_10,WX3590);
  and AND2_1025(WX2920,WX5038,WX2921);
  and AND2_1026(WX2923,WX3113,WX3590);
  and AND2_1027(WX2924,WX3745,WX2925);
  and AND2_1028(WX2929,WX2940,WX3589);
  and AND2_1029(WX2930,WX2936,WX2931);
  and AND2_1030(WX2933,CRC_OUT_7_9,WX3590);
  and AND2_1031(WX2934,WX5045,WX2935);
  and AND2_1032(WX2937,WX3115,WX3590);
  and AND2_1033(WX2938,WX3752,WX2939);
  and AND2_1034(WX2943,WX2954,WX3589);
  and AND2_1035(WX2944,WX2950,WX2945);
  and AND2_1036(WX2947,CRC_OUT_7_8,WX3590);
  and AND2_1037(WX2948,WX5052,WX2949);
  and AND2_1038(WX2951,WX3117,WX3590);
  and AND2_1039(WX2952,WX3759,WX2953);
  and AND2_1040(WX2957,WX2968,WX3589);
  and AND2_1041(WX2958,WX2964,WX2959);
  and AND2_1042(WX2961,CRC_OUT_7_7,WX3590);
  and AND2_1043(WX2962,WX5059,WX2963);
  and AND2_1044(WX2965,WX3119,WX3590);
  and AND2_1045(WX2966,WX3766,WX2967);
  and AND2_1046(WX2971,WX2982,WX3589);
  and AND2_1047(WX2972,WX2978,WX2973);
  and AND2_1048(WX2975,CRC_OUT_7_6,WX3590);
  and AND2_1049(WX2976,WX5066,WX2977);
  and AND2_1050(WX2979,WX3121,WX3590);
  and AND2_1051(WX2980,WX3773,WX2981);
  and AND2_1052(WX2985,WX2996,WX3589);
  and AND2_1053(WX2986,WX2992,WX2987);
  and AND2_1054(WX2989,CRC_OUT_7_5,WX3590);
  and AND2_1055(WX2990,WX5073,WX2991);
  and AND2_1056(WX2993,WX3123,WX3590);
  and AND2_1057(WX2994,WX3780,WX2995);
  and AND2_1058(WX2999,WX3010,WX3589);
  and AND2_1059(WX3000,WX3006,WX3001);
  and AND2_1060(WX3003,CRC_OUT_7_4,WX3590);
  and AND2_1061(WX3004,WX5080,WX3005);
  and AND2_1062(WX3007,WX3125,WX3590);
  and AND2_1063(WX3008,WX3787,WX3009);
  and AND2_1064(WX3013,WX3024,WX3589);
  and AND2_1065(WX3014,WX3020,WX3015);
  and AND2_1066(WX3017,CRC_OUT_7_3,WX3590);
  and AND2_1067(WX3018,WX5087,WX3019);
  and AND2_1068(WX3021,WX3127,WX3590);
  and AND2_1069(WX3022,WX3794,WX3023);
  and AND2_1070(WX3027,WX3038,WX3589);
  and AND2_1071(WX3028,WX3034,WX3029);
  and AND2_1072(WX3031,CRC_OUT_7_2,WX3590);
  and AND2_1073(WX3032,WX5094,WX3033);
  and AND2_1074(WX3035,WX3129,WX3590);
  and AND2_1075(WX3036,WX3801,WX3037);
  and AND2_1076(WX3041,WX3052,WX3589);
  and AND2_1077(WX3042,WX3048,WX3043);
  and AND2_1078(WX3045,CRC_OUT_7_1,WX3590);
  and AND2_1079(WX3046,WX5101,WX3047);
  and AND2_1080(WX3049,WX3131,WX3590);
  and AND2_1081(WX3050,WX3808,WX3051);
  and AND2_1082(WX3055,WX3066,WX3589);
  and AND2_1083(WX3056,WX3062,WX3057);
  and AND2_1084(WX3059,CRC_OUT_7_0,WX3590);
  and AND2_1085(WX3060,WX5108,WX3061);
  and AND2_1086(WX3063,WX3133,WX3590);
  and AND2_1087(WX3064,WX3815,WX3065);
  and AND2_1088(WX3070,WX3073,RESET);
  and AND2_1089(WX3072,WX3075,RESET);
  and AND2_1090(WX3074,WX3077,RESET);
  and AND2_1091(WX3076,WX3079,RESET);
  and AND2_1092(WX3078,WX3081,RESET);
  and AND2_1093(WX3080,WX3083,RESET);
  and AND2_1094(WX3082,WX3085,RESET);
  and AND2_1095(WX3084,WX3087,RESET);
  and AND2_1096(WX3086,WX3089,RESET);
  and AND2_1097(WX3088,WX3091,RESET);
  and AND2_1098(WX3090,WX3093,RESET);
  and AND2_1099(WX3092,WX3095,RESET);
  and AND2_1100(WX3094,WX3097,RESET);
  and AND2_1101(WX3096,WX3099,RESET);
  and AND2_1102(WX3098,WX3101,RESET);
  and AND2_1103(WX3100,WX3103,RESET);
  and AND2_1104(WX3102,WX3105,RESET);
  and AND2_1105(WX3104,WX3107,RESET);
  and AND2_1106(WX3106,WX3109,RESET);
  and AND2_1107(WX3108,WX3111,RESET);
  and AND2_1108(WX3110,WX3113,RESET);
  and AND2_1109(WX3112,WX3115,RESET);
  and AND2_1110(WX3114,WX3117,RESET);
  and AND2_1111(WX3116,WX3119,RESET);
  and AND2_1112(WX3118,WX3121,RESET);
  and AND2_1113(WX3120,WX3123,RESET);
  and AND2_1114(WX3122,WX3125,RESET);
  and AND2_1115(WX3124,WX3127,RESET);
  and AND2_1116(WX3126,WX3129,RESET);
  and AND2_1117(WX3128,WX3131,RESET);
  and AND2_1118(WX3130,WX3133,RESET);
  and AND2_1119(WX3132,WX3069,RESET);
  and AND2_1120(WX3230,WX2634,RESET);
  and AND2_1121(WX3232,WX2648,RESET);
  and AND2_1122(WX3234,WX2662,RESET);
  and AND2_1123(WX3236,WX2676,RESET);
  and AND2_1124(WX3238,WX2690,RESET);
  and AND2_1125(WX3240,WX2704,RESET);
  and AND2_1126(WX3242,WX2718,RESET);
  and AND2_1127(WX3244,WX2732,RESET);
  and AND2_1128(WX3246,WX2746,RESET);
  and AND2_1129(WX3248,WX2760,RESET);
  and AND2_1130(WX3250,WX2774,RESET);
  and AND2_1131(WX3252,WX2788,RESET);
  and AND2_1132(WX3254,WX2802,RESET);
  and AND2_1133(WX3256,WX2816,RESET);
  and AND2_1134(WX3258,WX2830,RESET);
  and AND2_1135(WX3260,WX2844,RESET);
  and AND2_1136(WX3262,WX2858,RESET);
  and AND2_1137(WX3264,WX2872,RESET);
  and AND2_1138(WX3266,WX2886,RESET);
  and AND2_1139(WX3268,WX2900,RESET);
  and AND2_1140(WX3270,WX2914,RESET);
  and AND2_1141(WX3272,WX2928,RESET);
  and AND2_1142(WX3274,WX2942,RESET);
  and AND2_1143(WX3276,WX2956,RESET);
  and AND2_1144(WX3278,WX2970,RESET);
  and AND2_1145(WX3280,WX2984,RESET);
  and AND2_1146(WX3282,WX2998,RESET);
  and AND2_1147(WX3284,WX3012,RESET);
  and AND2_1148(WX3286,WX3026,RESET);
  and AND2_1149(WX3288,WX3040,RESET);
  and AND2_1150(WX3290,WX3054,RESET);
  and AND2_1151(WX3292,WX3068,RESET);
  and AND2_1152(WX3294,WX3231,RESET);
  and AND2_1153(WX3296,WX3233,RESET);
  and AND2_1154(WX3298,WX3235,RESET);
  and AND2_1155(WX3300,WX3237,RESET);
  and AND2_1156(WX3302,WX3239,RESET);
  and AND2_1157(WX3304,WX3241,RESET);
  and AND2_1158(WX3306,WX3243,RESET);
  and AND2_1159(WX3308,WX3245,RESET);
  and AND2_1160(WX3310,WX3247,RESET);
  and AND2_1161(WX3312,WX3249,RESET);
  and AND2_1162(WX3314,WX3251,RESET);
  and AND2_1163(WX3316,WX3253,RESET);
  and AND2_1164(WX3318,WX3255,RESET);
  and AND2_1165(WX3320,WX3257,RESET);
  and AND2_1166(WX3322,WX3259,RESET);
  and AND2_1167(WX3324,WX3261,RESET);
  and AND2_1168(WX3326,WX3263,RESET);
  and AND2_1169(WX3328,WX3265,RESET);
  and AND2_1170(WX3330,WX3267,RESET);
  and AND2_1171(WX3332,WX3269,RESET);
  and AND2_1172(WX3334,WX3271,RESET);
  and AND2_1173(WX3336,WX3273,RESET);
  and AND2_1174(WX3338,WX3275,RESET);
  and AND2_1175(WX3340,WX3277,RESET);
  and AND2_1176(WX3342,WX3279,RESET);
  and AND2_1177(WX3344,WX3281,RESET);
  and AND2_1178(WX3346,WX3283,RESET);
  and AND2_1179(WX3348,WX3285,RESET);
  and AND2_1180(WX3350,WX3287,RESET);
  and AND2_1181(WX3352,WX3289,RESET);
  and AND2_1182(WX3354,WX3291,RESET);
  and AND2_1183(WX3356,WX3293,RESET);
  and AND2_1184(WX3358,WX3295,RESET);
  and AND2_1185(WX3360,WX3297,RESET);
  and AND2_1186(WX3362,WX3299,RESET);
  and AND2_1187(WX3364,WX3301,RESET);
  and AND2_1188(WX3366,WX3303,RESET);
  and AND2_1189(WX3368,WX3305,RESET);
  and AND2_1190(WX3370,WX3307,RESET);
  and AND2_1191(WX3372,WX3309,RESET);
  and AND2_1192(WX3374,WX3311,RESET);
  and AND2_1193(WX3376,WX3313,RESET);
  and AND2_1194(WX3378,WX3315,RESET);
  and AND2_1195(WX3380,WX3317,RESET);
  and AND2_1196(WX3382,WX3319,RESET);
  and AND2_1197(WX3384,WX3321,RESET);
  and AND2_1198(WX3386,WX3323,RESET);
  and AND2_1199(WX3388,WX3325,RESET);
  and AND2_1200(WX3390,WX3327,RESET);
  and AND2_1201(WX3392,WX3329,RESET);
  and AND2_1202(WX3394,WX3331,RESET);
  and AND2_1203(WX3396,WX3333,RESET);
  and AND2_1204(WX3398,WX3335,RESET);
  and AND2_1205(WX3400,WX3337,RESET);
  and AND2_1206(WX3402,WX3339,RESET);
  and AND2_1207(WX3404,WX3341,RESET);
  and AND2_1208(WX3406,WX3343,RESET);
  and AND2_1209(WX3408,WX3345,RESET);
  and AND2_1210(WX3410,WX3347,RESET);
  and AND2_1211(WX3412,WX3349,RESET);
  and AND2_1212(WX3414,WX3351,RESET);
  and AND2_1213(WX3416,WX3353,RESET);
  and AND2_1214(WX3418,WX3355,RESET);
  and AND2_1215(WX3420,WX3357,RESET);
  and AND2_1216(WX3422,WX3359,RESET);
  and AND2_1217(WX3424,WX3361,RESET);
  and AND2_1218(WX3426,WX3363,RESET);
  and AND2_1219(WX3428,WX3365,RESET);
  and AND2_1220(WX3430,WX3367,RESET);
  and AND2_1221(WX3432,WX3369,RESET);
  and AND2_1222(WX3434,WX3371,RESET);
  and AND2_1223(WX3436,WX3373,RESET);
  and AND2_1224(WX3438,WX3375,RESET);
  and AND2_1225(WX3440,WX3377,RESET);
  and AND2_1226(WX3442,WX3379,RESET);
  and AND2_1227(WX3444,WX3381,RESET);
  and AND2_1228(WX3446,WX3383,RESET);
  and AND2_1229(WX3448,WX3385,RESET);
  and AND2_1230(WX3450,WX3387,RESET);
  and AND2_1231(WX3452,WX3389,RESET);
  and AND2_1232(WX3454,WX3391,RESET);
  and AND2_1233(WX3456,WX3393,RESET);
  and AND2_1234(WX3458,WX3395,RESET);
  and AND2_1235(WX3460,WX3397,RESET);
  and AND2_1236(WX3462,WX3399,RESET);
  and AND2_1237(WX3464,WX3401,RESET);
  and AND2_1238(WX3466,WX3403,RESET);
  and AND2_1239(WX3468,WX3405,RESET);
  and AND2_1240(WX3470,WX3407,RESET);
  and AND2_1241(WX3472,WX3409,RESET);
  and AND2_1242(WX3474,WX3411,RESET);
  and AND2_1243(WX3476,WX3413,RESET);
  and AND2_1244(WX3478,WX3415,RESET);
  and AND2_1245(WX3480,WX3417,RESET);
  and AND2_1246(WX3482,WX3419,RESET);
  and AND2_1247(WX3484,WX3421,RESET);
  and AND2_1248(WX3593,WX3592,WX3591);
  and AND2_1249(WX3594,WX3166,WX3595);
  and AND2_1250(WX3600,WX3599,WX3591);
  and AND2_1251(WX3601,WX3167,WX3602);
  and AND2_1252(WX3607,WX3606,WX3591);
  and AND2_1253(WX3608,WX3168,WX3609);
  and AND2_1254(WX3614,WX3613,WX3591);
  and AND2_1255(WX3615,WX3169,WX3616);
  and AND2_1256(WX3621,WX3620,WX3591);
  and AND2_1257(WX3622,WX3170,WX3623);
  and AND2_1258(WX3628,WX3627,WX3591);
  and AND2_1259(WX3629,WX3171,WX3630);
  and AND2_1260(WX3635,WX3634,WX3591);
  and AND2_1261(WX3636,WX3172,WX3637);
  and AND2_1262(WX3642,WX3641,WX3591);
  and AND2_1263(WX3643,WX3173,WX3644);
  and AND2_1264(WX3649,WX3648,WX3591);
  and AND2_1265(WX3650,WX3174,WX3651);
  and AND2_1266(WX3656,WX3655,WX3591);
  and AND2_1267(WX3657,WX3175,WX3658);
  and AND2_1268(WX3663,WX3662,WX3591);
  and AND2_1269(WX3664,WX3176,WX3665);
  and AND2_1270(WX3670,WX3669,WX3591);
  and AND2_1271(WX3671,WX3177,WX3672);
  and AND2_1272(WX3677,WX3676,WX3591);
  and AND2_1273(WX3678,WX3178,WX3679);
  and AND2_1274(WX3684,WX3683,WX3591);
  and AND2_1275(WX3685,WX3179,WX3686);
  and AND2_1276(WX3691,WX3690,WX3591);
  and AND2_1277(WX3692,WX3180,WX3693);
  and AND2_1278(WX3698,WX3697,WX3591);
  and AND2_1279(WX3699,WX3181,WX3700);
  and AND2_1280(WX3705,WX3704,WX3591);
  and AND2_1281(WX3706,WX3182,WX3707);
  and AND2_1282(WX3712,WX3711,WX3591);
  and AND2_1283(WX3713,WX3183,WX3714);
  and AND2_1284(WX3719,WX3718,WX3591);
  and AND2_1285(WX3720,WX3184,WX3721);
  and AND2_1286(WX3726,WX3725,WX3591);
  and AND2_1287(WX3727,WX3185,WX3728);
  and AND2_1288(WX3733,WX3732,WX3591);
  and AND2_1289(WX3734,WX3186,WX3735);
  and AND2_1290(WX3740,WX3739,WX3591);
  and AND2_1291(WX3741,WX3187,WX3742);
  and AND2_1292(WX3747,WX3746,WX3591);
  and AND2_1293(WX3748,WX3188,WX3749);
  and AND2_1294(WX3754,WX3753,WX3591);
  and AND2_1295(WX3755,WX3189,WX3756);
  and AND2_1296(WX3761,WX3760,WX3591);
  and AND2_1297(WX3762,WX3190,WX3763);
  and AND2_1298(WX3768,WX3767,WX3591);
  and AND2_1299(WX3769,WX3191,WX3770);
  and AND2_1300(WX3775,WX3774,WX3591);
  and AND2_1301(WX3776,WX3192,WX3777);
  and AND2_1302(WX3782,WX3781,WX3591);
  and AND2_1303(WX3783,WX3193,WX3784);
  and AND2_1304(WX3789,WX3788,WX3591);
  and AND2_1305(WX3790,WX3194,WX3791);
  and AND2_1306(WX3796,WX3795,WX3591);
  and AND2_1307(WX3797,WX3195,WX3798);
  and AND2_1308(WX3803,WX3802,WX3591);
  and AND2_1309(WX3804,WX3196,WX3805);
  and AND2_1310(WX3810,WX3809,WX3591);
  and AND2_1311(WX3811,WX3197,WX3812);
  and AND2_1312(WX3850,WX3820,WX3849);
  and AND2_1313(WX3852,WX3848,WX3849);
  and AND2_1314(WX3854,WX3847,WX3849);
  and AND2_1315(WX3856,WX3846,WX3849);
  and AND2_1316(WX3858,WX3819,WX3849);
  and AND2_1317(WX3860,WX3845,WX3849);
  and AND2_1318(WX3862,WX3844,WX3849);
  and AND2_1319(WX3864,WX3843,WX3849);
  and AND2_1320(WX3866,WX3842,WX3849);
  and AND2_1321(WX3868,WX3841,WX3849);
  and AND2_1322(WX3870,WX3840,WX3849);
  and AND2_1323(WX3872,WX3818,WX3849);
  and AND2_1324(WX3874,WX3839,WX3849);
  and AND2_1325(WX3876,WX3838,WX3849);
  and AND2_1326(WX3878,WX3837,WX3849);
  and AND2_1327(WX3880,WX3836,WX3849);
  and AND2_1328(WX3882,WX3817,WX3849);
  and AND2_1329(WX3884,WX3835,WX3849);
  and AND2_1330(WX3886,WX3834,WX3849);
  and AND2_1331(WX3888,WX3833,WX3849);
  and AND2_1332(WX3890,WX3832,WX3849);
  and AND2_1333(WX3892,WX3831,WX3849);
  and AND2_1334(WX3894,WX3830,WX3849);
  and AND2_1335(WX3896,WX3829,WX3849);
  and AND2_1336(WX3898,WX3828,WX3849);
  and AND2_1337(WX3900,WX3827,WX3849);
  and AND2_1338(WX3902,WX3826,WX3849);
  and AND2_1339(WX3904,WX3825,WX3849);
  and AND2_1340(WX3906,WX3824,WX3849);
  and AND2_1341(WX3908,WX3823,WX3849);
  and AND2_1342(WX3910,WX3822,WX3849);
  and AND2_1343(WX3912,WX3821,WX3849);
  and AND2_1344(WX3914,WX3925,WX4882);
  and AND2_1345(WX3915,WX3921,WX3916);
  and AND2_1346(WX3918,CRC_OUT_6_31,WX4883);
  and AND2_1347(WX3919,WX6184,WX3920);
  and AND2_1348(WX3922,WX4364,WX4883);
  and AND2_1349(WX3923,WX4891,WX3924);
  and AND2_1350(WX3928,WX3939,WX4882);
  and AND2_1351(WX3929,WX3935,WX3930);
  and AND2_1352(WX3932,CRC_OUT_6_30,WX4883);
  and AND2_1353(WX3933,WX6191,WX3934);
  and AND2_1354(WX3936,WX4366,WX4883);
  and AND2_1355(WX3937,WX4898,WX3938);
  and AND2_1356(WX3942,WX3953,WX4882);
  and AND2_1357(WX3943,WX3949,WX3944);
  and AND2_1358(WX3946,CRC_OUT_6_29,WX4883);
  and AND2_1359(WX3947,WX6198,WX3948);
  and AND2_1360(WX3950,WX4368,WX4883);
  and AND2_1361(WX3951,WX4905,WX3952);
  and AND2_1362(WX3956,WX3967,WX4882);
  and AND2_1363(WX3957,WX3963,WX3958);
  and AND2_1364(WX3960,CRC_OUT_6_28,WX4883);
  and AND2_1365(WX3961,WX6205,WX3962);
  and AND2_1366(WX3964,WX4370,WX4883);
  and AND2_1367(WX3965,WX4912,WX3966);
  and AND2_1368(WX3970,WX3981,WX4882);
  and AND2_1369(WX3971,WX3977,WX3972);
  and AND2_1370(WX3974,CRC_OUT_6_27,WX4883);
  and AND2_1371(WX3975,WX6212,WX3976);
  and AND2_1372(WX3978,WX4372,WX4883);
  and AND2_1373(WX3979,WX4919,WX3980);
  and AND2_1374(WX3984,WX3995,WX4882);
  and AND2_1375(WX3985,WX3991,WX3986);
  and AND2_1376(WX3988,CRC_OUT_6_26,WX4883);
  and AND2_1377(WX3989,WX6219,WX3990);
  and AND2_1378(WX3992,WX4374,WX4883);
  and AND2_1379(WX3993,WX4926,WX3994);
  and AND2_1380(WX3998,WX4009,WX4882);
  and AND2_1381(WX3999,WX4005,WX4000);
  and AND2_1382(WX4002,CRC_OUT_6_25,WX4883);
  and AND2_1383(WX4003,WX6226,WX4004);
  and AND2_1384(WX4006,WX4376,WX4883);
  and AND2_1385(WX4007,WX4933,WX4008);
  and AND2_1386(WX4012,WX4023,WX4882);
  and AND2_1387(WX4013,WX4019,WX4014);
  and AND2_1388(WX4016,CRC_OUT_6_24,WX4883);
  and AND2_1389(WX4017,WX6233,WX4018);
  and AND2_1390(WX4020,WX4378,WX4883);
  and AND2_1391(WX4021,WX4940,WX4022);
  and AND2_1392(WX4026,WX4037,WX4882);
  and AND2_1393(WX4027,WX4033,WX4028);
  and AND2_1394(WX4030,CRC_OUT_6_23,WX4883);
  and AND2_1395(WX4031,WX6240,WX4032);
  and AND2_1396(WX4034,WX4380,WX4883);
  and AND2_1397(WX4035,WX4947,WX4036);
  and AND2_1398(WX4040,WX4051,WX4882);
  and AND2_1399(WX4041,WX4047,WX4042);
  and AND2_1400(WX4044,CRC_OUT_6_22,WX4883);
  and AND2_1401(WX4045,WX6247,WX4046);
  and AND2_1402(WX4048,WX4382,WX4883);
  and AND2_1403(WX4049,WX4954,WX4050);
  and AND2_1404(WX4054,WX4065,WX4882);
  and AND2_1405(WX4055,WX4061,WX4056);
  and AND2_1406(WX4058,CRC_OUT_6_21,WX4883);
  and AND2_1407(WX4059,WX6254,WX4060);
  and AND2_1408(WX4062,WX4384,WX4883);
  and AND2_1409(WX4063,WX4961,WX4064);
  and AND2_1410(WX4068,WX4079,WX4882);
  and AND2_1411(WX4069,WX4075,WX4070);
  and AND2_1412(WX4072,CRC_OUT_6_20,WX4883);
  and AND2_1413(WX4073,WX6261,WX4074);
  and AND2_1414(WX4076,WX4386,WX4883);
  and AND2_1415(WX4077,WX4968,WX4078);
  and AND2_1416(WX4082,WX4093,WX4882);
  and AND2_1417(WX4083,WX4089,WX4084);
  and AND2_1418(WX4086,CRC_OUT_6_19,WX4883);
  and AND2_1419(WX4087,WX6268,WX4088);
  and AND2_1420(WX4090,WX4388,WX4883);
  and AND2_1421(WX4091,WX4975,WX4092);
  and AND2_1422(WX4096,WX4107,WX4882);
  and AND2_1423(WX4097,WX4103,WX4098);
  and AND2_1424(WX4100,CRC_OUT_6_18,WX4883);
  and AND2_1425(WX4101,WX6275,WX4102);
  and AND2_1426(WX4104,WX4390,WX4883);
  and AND2_1427(WX4105,WX4982,WX4106);
  and AND2_1428(WX4110,WX4121,WX4882);
  and AND2_1429(WX4111,WX4117,WX4112);
  and AND2_1430(WX4114,CRC_OUT_6_17,WX4883);
  and AND2_1431(WX4115,WX6282,WX4116);
  and AND2_1432(WX4118,WX4392,WX4883);
  and AND2_1433(WX4119,WX4989,WX4120);
  and AND2_1434(WX4124,WX4135,WX4882);
  and AND2_1435(WX4125,WX4131,WX4126);
  and AND2_1436(WX4128,CRC_OUT_6_16,WX4883);
  and AND2_1437(WX4129,WX6289,WX4130);
  and AND2_1438(WX4132,WX4394,WX4883);
  and AND2_1439(WX4133,WX4996,WX4134);
  and AND2_1440(WX4138,WX4149,WX4882);
  and AND2_1441(WX4139,WX4145,WX4140);
  and AND2_1442(WX4142,CRC_OUT_6_15,WX4883);
  and AND2_1443(WX4143,WX6296,WX4144);
  and AND2_1444(WX4146,WX4396,WX4883);
  and AND2_1445(WX4147,WX5003,WX4148);
  and AND2_1446(WX4152,WX4163,WX4882);
  and AND2_1447(WX4153,WX4159,WX4154);
  and AND2_1448(WX4156,CRC_OUT_6_14,WX4883);
  and AND2_1449(WX4157,WX6303,WX4158);
  and AND2_1450(WX4160,WX4398,WX4883);
  and AND2_1451(WX4161,WX5010,WX4162);
  and AND2_1452(WX4166,WX4177,WX4882);
  and AND2_1453(WX4167,WX4173,WX4168);
  and AND2_1454(WX4170,CRC_OUT_6_13,WX4883);
  and AND2_1455(WX4171,WX6310,WX4172);
  and AND2_1456(WX4174,WX4400,WX4883);
  and AND2_1457(WX4175,WX5017,WX4176);
  and AND2_1458(WX4180,WX4191,WX4882);
  and AND2_1459(WX4181,WX4187,WX4182);
  and AND2_1460(WX4184,CRC_OUT_6_12,WX4883);
  and AND2_1461(WX4185,WX6317,WX4186);
  and AND2_1462(WX4188,WX4402,WX4883);
  and AND2_1463(WX4189,WX5024,WX4190);
  and AND2_1464(WX4194,WX4205,WX4882);
  and AND2_1465(WX4195,WX4201,WX4196);
  and AND2_1466(WX4198,CRC_OUT_6_11,WX4883);
  and AND2_1467(WX4199,WX6324,WX4200);
  and AND2_1468(WX4202,WX4404,WX4883);
  and AND2_1469(WX4203,WX5031,WX4204);
  and AND2_1470(WX4208,WX4219,WX4882);
  and AND2_1471(WX4209,WX4215,WX4210);
  and AND2_1472(WX4212,CRC_OUT_6_10,WX4883);
  and AND2_1473(WX4213,WX6331,WX4214);
  and AND2_1474(WX4216,WX4406,WX4883);
  and AND2_1475(WX4217,WX5038,WX4218);
  and AND2_1476(WX4222,WX4233,WX4882);
  and AND2_1477(WX4223,WX4229,WX4224);
  and AND2_1478(WX4226,CRC_OUT_6_9,WX4883);
  and AND2_1479(WX4227,WX6338,WX4228);
  and AND2_1480(WX4230,WX4408,WX4883);
  and AND2_1481(WX4231,WX5045,WX4232);
  and AND2_1482(WX4236,WX4247,WX4882);
  and AND2_1483(WX4237,WX4243,WX4238);
  and AND2_1484(WX4240,CRC_OUT_6_8,WX4883);
  and AND2_1485(WX4241,WX6345,WX4242);
  and AND2_1486(WX4244,WX4410,WX4883);
  and AND2_1487(WX4245,WX5052,WX4246);
  and AND2_1488(WX4250,WX4261,WX4882);
  and AND2_1489(WX4251,WX4257,WX4252);
  and AND2_1490(WX4254,CRC_OUT_6_7,WX4883);
  and AND2_1491(WX4255,WX6352,WX4256);
  and AND2_1492(WX4258,WX4412,WX4883);
  and AND2_1493(WX4259,WX5059,WX4260);
  and AND2_1494(WX4264,WX4275,WX4882);
  and AND2_1495(WX4265,WX4271,WX4266);
  and AND2_1496(WX4268,CRC_OUT_6_6,WX4883);
  and AND2_1497(WX4269,WX6359,WX4270);
  and AND2_1498(WX4272,WX4414,WX4883);
  and AND2_1499(WX4273,WX5066,WX4274);
  and AND2_1500(WX4278,WX4289,WX4882);
  and AND2_1501(WX4279,WX4285,WX4280);
  and AND2_1502(WX4282,CRC_OUT_6_5,WX4883);
  and AND2_1503(WX4283,WX6366,WX4284);
  and AND2_1504(WX4286,WX4416,WX4883);
  and AND2_1505(WX4287,WX5073,WX4288);
  and AND2_1506(WX4292,WX4303,WX4882);
  and AND2_1507(WX4293,WX4299,WX4294);
  and AND2_1508(WX4296,CRC_OUT_6_4,WX4883);
  and AND2_1509(WX4297,WX6373,WX4298);
  and AND2_1510(WX4300,WX4418,WX4883);
  and AND2_1511(WX4301,WX5080,WX4302);
  and AND2_1512(WX4306,WX4317,WX4882);
  and AND2_1513(WX4307,WX4313,WX4308);
  and AND2_1514(WX4310,CRC_OUT_6_3,WX4883);
  and AND2_1515(WX4311,WX6380,WX4312);
  and AND2_1516(WX4314,WX4420,WX4883);
  and AND2_1517(WX4315,WX5087,WX4316);
  and AND2_1518(WX4320,WX4331,WX4882);
  and AND2_1519(WX4321,WX4327,WX4322);
  and AND2_1520(WX4324,CRC_OUT_6_2,WX4883);
  and AND2_1521(WX4325,WX6387,WX4326);
  and AND2_1522(WX4328,WX4422,WX4883);
  and AND2_1523(WX4329,WX5094,WX4330);
  and AND2_1524(WX4334,WX4345,WX4882);
  and AND2_1525(WX4335,WX4341,WX4336);
  and AND2_1526(WX4338,CRC_OUT_6_1,WX4883);
  and AND2_1527(WX4339,WX6394,WX4340);
  and AND2_1528(WX4342,WX4424,WX4883);
  and AND2_1529(WX4343,WX5101,WX4344);
  and AND2_1530(WX4348,WX4359,WX4882);
  and AND2_1531(WX4349,WX4355,WX4350);
  and AND2_1532(WX4352,CRC_OUT_6_0,WX4883);
  and AND2_1533(WX4353,WX6401,WX4354);
  and AND2_1534(WX4356,WX4426,WX4883);
  and AND2_1535(WX4357,WX5108,WX4358);
  and AND2_1536(WX4363,WX4366,RESET);
  and AND2_1537(WX4365,WX4368,RESET);
  and AND2_1538(WX4367,WX4370,RESET);
  and AND2_1539(WX4369,WX4372,RESET);
  and AND2_1540(WX4371,WX4374,RESET);
  and AND2_1541(WX4373,WX4376,RESET);
  and AND2_1542(WX4375,WX4378,RESET);
  and AND2_1543(WX4377,WX4380,RESET);
  and AND2_1544(WX4379,WX4382,RESET);
  and AND2_1545(WX4381,WX4384,RESET);
  and AND2_1546(WX4383,WX4386,RESET);
  and AND2_1547(WX4385,WX4388,RESET);
  and AND2_1548(WX4387,WX4390,RESET);
  and AND2_1549(WX4389,WX4392,RESET);
  and AND2_1550(WX4391,WX4394,RESET);
  and AND2_1551(WX4393,WX4396,RESET);
  and AND2_1552(WX4395,WX4398,RESET);
  and AND2_1553(WX4397,WX4400,RESET);
  and AND2_1554(WX4399,WX4402,RESET);
  and AND2_1555(WX4401,WX4404,RESET);
  and AND2_1556(WX4403,WX4406,RESET);
  and AND2_1557(WX4405,WX4408,RESET);
  and AND2_1558(WX4407,WX4410,RESET);
  and AND2_1559(WX4409,WX4412,RESET);
  and AND2_1560(WX4411,WX4414,RESET);
  and AND2_1561(WX4413,WX4416,RESET);
  and AND2_1562(WX4415,WX4418,RESET);
  and AND2_1563(WX4417,WX4420,RESET);
  and AND2_1564(WX4419,WX4422,RESET);
  and AND2_1565(WX4421,WX4424,RESET);
  and AND2_1566(WX4423,WX4426,RESET);
  and AND2_1567(WX4425,WX4362,RESET);
  and AND2_1568(WX4523,WX3927,RESET);
  and AND2_1569(WX4525,WX3941,RESET);
  and AND2_1570(WX4527,WX3955,RESET);
  and AND2_1571(WX4529,WX3969,RESET);
  and AND2_1572(WX4531,WX3983,RESET);
  and AND2_1573(WX4533,WX3997,RESET);
  and AND2_1574(WX4535,WX4011,RESET);
  and AND2_1575(WX4537,WX4025,RESET);
  and AND2_1576(WX4539,WX4039,RESET);
  and AND2_1577(WX4541,WX4053,RESET);
  and AND2_1578(WX4543,WX4067,RESET);
  and AND2_1579(WX4545,WX4081,RESET);
  and AND2_1580(WX4547,WX4095,RESET);
  and AND2_1581(WX4549,WX4109,RESET);
  and AND2_1582(WX4551,WX4123,RESET);
  and AND2_1583(WX4553,WX4137,RESET);
  and AND2_1584(WX4555,WX4151,RESET);
  and AND2_1585(WX4557,WX4165,RESET);
  and AND2_1586(WX4559,WX4179,RESET);
  and AND2_1587(WX4561,WX4193,RESET);
  and AND2_1588(WX4563,WX4207,RESET);
  and AND2_1589(WX4565,WX4221,RESET);
  and AND2_1590(WX4567,WX4235,RESET);
  and AND2_1591(WX4569,WX4249,RESET);
  and AND2_1592(WX4571,WX4263,RESET);
  and AND2_1593(WX4573,WX4277,RESET);
  and AND2_1594(WX4575,WX4291,RESET);
  and AND2_1595(WX4577,WX4305,RESET);
  and AND2_1596(WX4579,WX4319,RESET);
  and AND2_1597(WX4581,WX4333,RESET);
  and AND2_1598(WX4583,WX4347,RESET);
  and AND2_1599(WX4585,WX4361,RESET);
  and AND2_1600(WX4587,WX4524,RESET);
  and AND2_1601(WX4589,WX4526,RESET);
  and AND2_1602(WX4591,WX4528,RESET);
  and AND2_1603(WX4593,WX4530,RESET);
  and AND2_1604(WX4595,WX4532,RESET);
  and AND2_1605(WX4597,WX4534,RESET);
  and AND2_1606(WX4599,WX4536,RESET);
  and AND2_1607(WX4601,WX4538,RESET);
  and AND2_1608(WX4603,WX4540,RESET);
  and AND2_1609(WX4605,WX4542,RESET);
  and AND2_1610(WX4607,WX4544,RESET);
  and AND2_1611(WX4609,WX4546,RESET);
  and AND2_1612(WX4611,WX4548,RESET);
  and AND2_1613(WX4613,WX4550,RESET);
  and AND2_1614(WX4615,WX4552,RESET);
  and AND2_1615(WX4617,WX4554,RESET);
  and AND2_1616(WX4619,WX4556,RESET);
  and AND2_1617(WX4621,WX4558,RESET);
  and AND2_1618(WX4623,WX4560,RESET);
  and AND2_1619(WX4625,WX4562,RESET);
  and AND2_1620(WX4627,WX4564,RESET);
  and AND2_1621(WX4629,WX4566,RESET);
  and AND2_1622(WX4631,WX4568,RESET);
  and AND2_1623(WX4633,WX4570,RESET);
  and AND2_1624(WX4635,WX4572,RESET);
  and AND2_1625(WX4637,WX4574,RESET);
  and AND2_1626(WX4639,WX4576,RESET);
  and AND2_1627(WX4641,WX4578,RESET);
  and AND2_1628(WX4643,WX4580,RESET);
  and AND2_1629(WX4645,WX4582,RESET);
  and AND2_1630(WX4647,WX4584,RESET);
  and AND2_1631(WX4649,WX4586,RESET);
  and AND2_1632(WX4651,WX4588,RESET);
  and AND2_1633(WX4653,WX4590,RESET);
  and AND2_1634(WX4655,WX4592,RESET);
  and AND2_1635(WX4657,WX4594,RESET);
  and AND2_1636(WX4659,WX4596,RESET);
  and AND2_1637(WX4661,WX4598,RESET);
  and AND2_1638(WX4663,WX4600,RESET);
  and AND2_1639(WX4665,WX4602,RESET);
  and AND2_1640(WX4667,WX4604,RESET);
  and AND2_1641(WX4669,WX4606,RESET);
  and AND2_1642(WX4671,WX4608,RESET);
  and AND2_1643(WX4673,WX4610,RESET);
  and AND2_1644(WX4675,WX4612,RESET);
  and AND2_1645(WX4677,WX4614,RESET);
  and AND2_1646(WX4679,WX4616,RESET);
  and AND2_1647(WX4681,WX4618,RESET);
  and AND2_1648(WX4683,WX4620,RESET);
  and AND2_1649(WX4685,WX4622,RESET);
  and AND2_1650(WX4687,WX4624,RESET);
  and AND2_1651(WX4689,WX4626,RESET);
  and AND2_1652(WX4691,WX4628,RESET);
  and AND2_1653(WX4693,WX4630,RESET);
  and AND2_1654(WX4695,WX4632,RESET);
  and AND2_1655(WX4697,WX4634,RESET);
  and AND2_1656(WX4699,WX4636,RESET);
  and AND2_1657(WX4701,WX4638,RESET);
  and AND2_1658(WX4703,WX4640,RESET);
  and AND2_1659(WX4705,WX4642,RESET);
  and AND2_1660(WX4707,WX4644,RESET);
  and AND2_1661(WX4709,WX4646,RESET);
  and AND2_1662(WX4711,WX4648,RESET);
  and AND2_1663(WX4713,WX4650,RESET);
  and AND2_1664(WX4715,WX4652,RESET);
  and AND2_1665(WX4717,WX4654,RESET);
  and AND2_1666(WX4719,WX4656,RESET);
  and AND2_1667(WX4721,WX4658,RESET);
  and AND2_1668(WX4723,WX4660,RESET);
  and AND2_1669(WX4725,WX4662,RESET);
  and AND2_1670(WX4727,WX4664,RESET);
  and AND2_1671(WX4729,WX4666,RESET);
  and AND2_1672(WX4731,WX4668,RESET);
  and AND2_1673(WX4733,WX4670,RESET);
  and AND2_1674(WX4735,WX4672,RESET);
  and AND2_1675(WX4737,WX4674,RESET);
  and AND2_1676(WX4739,WX4676,RESET);
  and AND2_1677(WX4741,WX4678,RESET);
  and AND2_1678(WX4743,WX4680,RESET);
  and AND2_1679(WX4745,WX4682,RESET);
  and AND2_1680(WX4747,WX4684,RESET);
  and AND2_1681(WX4749,WX4686,RESET);
  and AND2_1682(WX4751,WX4688,RESET);
  and AND2_1683(WX4753,WX4690,RESET);
  and AND2_1684(WX4755,WX4692,RESET);
  and AND2_1685(WX4757,WX4694,RESET);
  and AND2_1686(WX4759,WX4696,RESET);
  and AND2_1687(WX4761,WX4698,RESET);
  and AND2_1688(WX4763,WX4700,RESET);
  and AND2_1689(WX4765,WX4702,RESET);
  and AND2_1690(WX4767,WX4704,RESET);
  and AND2_1691(WX4769,WX4706,RESET);
  and AND2_1692(WX4771,WX4708,RESET);
  and AND2_1693(WX4773,WX4710,RESET);
  and AND2_1694(WX4775,WX4712,RESET);
  and AND2_1695(WX4777,WX4714,RESET);
  and AND2_1696(WX4886,WX4885,WX4884);
  and AND2_1697(WX4887,WX4459,WX4888);
  and AND2_1698(WX4893,WX4892,WX4884);
  and AND2_1699(WX4894,WX4460,WX4895);
  and AND2_1700(WX4900,WX4899,WX4884);
  and AND2_1701(WX4901,WX4461,WX4902);
  and AND2_1702(WX4907,WX4906,WX4884);
  and AND2_1703(WX4908,WX4462,WX4909);
  and AND2_1704(WX4914,WX4913,WX4884);
  and AND2_1705(WX4915,WX4463,WX4916);
  and AND2_1706(WX4921,WX4920,WX4884);
  and AND2_1707(WX4922,WX4464,WX4923);
  and AND2_1708(WX4928,WX4927,WX4884);
  and AND2_1709(WX4929,WX4465,WX4930);
  and AND2_1710(WX4935,WX4934,WX4884);
  and AND2_1711(WX4936,WX4466,WX4937);
  and AND2_1712(WX4942,WX4941,WX4884);
  and AND2_1713(WX4943,WX4467,WX4944);
  and AND2_1714(WX4949,WX4948,WX4884);
  and AND2_1715(WX4950,WX4468,WX4951);
  and AND2_1716(WX4956,WX4955,WX4884);
  and AND2_1717(WX4957,WX4469,WX4958);
  and AND2_1718(WX4963,WX4962,WX4884);
  and AND2_1719(WX4964,WX4470,WX4965);
  and AND2_1720(WX4970,WX4969,WX4884);
  and AND2_1721(WX4971,WX4471,WX4972);
  and AND2_1722(WX4977,WX4976,WX4884);
  and AND2_1723(WX4978,WX4472,WX4979);
  and AND2_1724(WX4984,WX4983,WX4884);
  and AND2_1725(WX4985,WX4473,WX4986);
  and AND2_1726(WX4991,WX4990,WX4884);
  and AND2_1727(WX4992,WX4474,WX4993);
  and AND2_1728(WX4998,WX4997,WX4884);
  and AND2_1729(WX4999,WX4475,WX5000);
  and AND2_1730(WX5005,WX5004,WX4884);
  and AND2_1731(WX5006,WX4476,WX5007);
  and AND2_1732(WX5012,WX5011,WX4884);
  and AND2_1733(WX5013,WX4477,WX5014);
  and AND2_1734(WX5019,WX5018,WX4884);
  and AND2_1735(WX5020,WX4478,WX5021);
  and AND2_1736(WX5026,WX5025,WX4884);
  and AND2_1737(WX5027,WX4479,WX5028);
  and AND2_1738(WX5033,WX5032,WX4884);
  and AND2_1739(WX5034,WX4480,WX5035);
  and AND2_1740(WX5040,WX5039,WX4884);
  and AND2_1741(WX5041,WX4481,WX5042);
  and AND2_1742(WX5047,WX5046,WX4884);
  and AND2_1743(WX5048,WX4482,WX5049);
  and AND2_1744(WX5054,WX5053,WX4884);
  and AND2_1745(WX5055,WX4483,WX5056);
  and AND2_1746(WX5061,WX5060,WX4884);
  and AND2_1747(WX5062,WX4484,WX5063);
  and AND2_1748(WX5068,WX5067,WX4884);
  and AND2_1749(WX5069,WX4485,WX5070);
  and AND2_1750(WX5075,WX5074,WX4884);
  and AND2_1751(WX5076,WX4486,WX5077);
  and AND2_1752(WX5082,WX5081,WX4884);
  and AND2_1753(WX5083,WX4487,WX5084);
  and AND2_1754(WX5089,WX5088,WX4884);
  and AND2_1755(WX5090,WX4488,WX5091);
  and AND2_1756(WX5096,WX5095,WX4884);
  and AND2_1757(WX5097,WX4489,WX5098);
  and AND2_1758(WX5103,WX5102,WX4884);
  and AND2_1759(WX5104,WX4490,WX5105);
  and AND2_1760(WX5143,WX5113,WX5142);
  and AND2_1761(WX5145,WX5141,WX5142);
  and AND2_1762(WX5147,WX5140,WX5142);
  and AND2_1763(WX5149,WX5139,WX5142);
  and AND2_1764(WX5151,WX5112,WX5142);
  and AND2_1765(WX5153,WX5138,WX5142);
  and AND2_1766(WX5155,WX5137,WX5142);
  and AND2_1767(WX5157,WX5136,WX5142);
  and AND2_1768(WX5159,WX5135,WX5142);
  and AND2_1769(WX5161,WX5134,WX5142);
  and AND2_1770(WX5163,WX5133,WX5142);
  and AND2_1771(WX5165,WX5111,WX5142);
  and AND2_1772(WX5167,WX5132,WX5142);
  and AND2_1773(WX5169,WX5131,WX5142);
  and AND2_1774(WX5171,WX5130,WX5142);
  and AND2_1775(WX5173,WX5129,WX5142);
  and AND2_1776(WX5175,WX5110,WX5142);
  and AND2_1777(WX5177,WX5128,WX5142);
  and AND2_1778(WX5179,WX5127,WX5142);
  and AND2_1779(WX5181,WX5126,WX5142);
  and AND2_1780(WX5183,WX5125,WX5142);
  and AND2_1781(WX5185,WX5124,WX5142);
  and AND2_1782(WX5187,WX5123,WX5142);
  and AND2_1783(WX5189,WX5122,WX5142);
  and AND2_1784(WX5191,WX5121,WX5142);
  and AND2_1785(WX5193,WX5120,WX5142);
  and AND2_1786(WX5195,WX5119,WX5142);
  and AND2_1787(WX5197,WX5118,WX5142);
  and AND2_1788(WX5199,WX5117,WX5142);
  and AND2_1789(WX5201,WX5116,WX5142);
  and AND2_1790(WX5203,WX5115,WX5142);
  and AND2_1791(WX5205,WX5114,WX5142);
  and AND2_1792(WX5207,WX5218,WX6175);
  and AND2_1793(WX5208,WX5214,WX5209);
  and AND2_1794(WX5211,CRC_OUT_5_31,WX6176);
  and AND2_1795(WX5212,WX7477,WX5213);
  and AND2_1796(WX5215,WX5657,WX6176);
  and AND2_1797(WX5216,WX6184,WX5217);
  and AND2_1798(WX5221,WX5232,WX6175);
  and AND2_1799(WX5222,WX5228,WX5223);
  and AND2_1800(WX5225,CRC_OUT_5_30,WX6176);
  and AND2_1801(WX5226,WX7484,WX5227);
  and AND2_1802(WX5229,WX5659,WX6176);
  and AND2_1803(WX5230,WX6191,WX5231);
  and AND2_1804(WX5235,WX5246,WX6175);
  and AND2_1805(WX5236,WX5242,WX5237);
  and AND2_1806(WX5239,CRC_OUT_5_29,WX6176);
  and AND2_1807(WX5240,WX7491,WX5241);
  and AND2_1808(WX5243,WX5661,WX6176);
  and AND2_1809(WX5244,WX6198,WX5245);
  and AND2_1810(WX5249,WX5260,WX6175);
  and AND2_1811(WX5250,WX5256,WX5251);
  and AND2_1812(WX5253,CRC_OUT_5_28,WX6176);
  and AND2_1813(WX5254,WX7498,WX5255);
  and AND2_1814(WX5257,WX5663,WX6176);
  and AND2_1815(WX5258,WX6205,WX5259);
  and AND2_1816(WX5263,WX5274,WX6175);
  and AND2_1817(WX5264,WX5270,WX5265);
  and AND2_1818(WX5267,CRC_OUT_5_27,WX6176);
  and AND2_1819(WX5268,WX7505,WX5269);
  and AND2_1820(WX5271,WX5665,WX6176);
  and AND2_1821(WX5272,WX6212,WX5273);
  and AND2_1822(WX5277,WX5288,WX6175);
  and AND2_1823(WX5278,WX5284,WX5279);
  and AND2_1824(WX5281,CRC_OUT_5_26,WX6176);
  and AND2_1825(WX5282,WX7512,WX5283);
  and AND2_1826(WX5285,WX5667,WX6176);
  and AND2_1827(WX5286,WX6219,WX5287);
  and AND2_1828(WX5291,WX5302,WX6175);
  and AND2_1829(WX5292,WX5298,WX5293);
  and AND2_1830(WX5295,CRC_OUT_5_25,WX6176);
  and AND2_1831(WX5296,WX7519,WX5297);
  and AND2_1832(WX5299,WX5669,WX6176);
  and AND2_1833(WX5300,WX6226,WX5301);
  and AND2_1834(WX5305,WX5316,WX6175);
  and AND2_1835(WX5306,WX5312,WX5307);
  and AND2_1836(WX5309,CRC_OUT_5_24,WX6176);
  and AND2_1837(WX5310,WX7526,WX5311);
  and AND2_1838(WX5313,WX5671,WX6176);
  and AND2_1839(WX5314,WX6233,WX5315);
  and AND2_1840(WX5319,WX5330,WX6175);
  and AND2_1841(WX5320,WX5326,WX5321);
  and AND2_1842(WX5323,CRC_OUT_5_23,WX6176);
  and AND2_1843(WX5324,WX7533,WX5325);
  and AND2_1844(WX5327,WX5673,WX6176);
  and AND2_1845(WX5328,WX6240,WX5329);
  and AND2_1846(WX5333,WX5344,WX6175);
  and AND2_1847(WX5334,WX5340,WX5335);
  and AND2_1848(WX5337,CRC_OUT_5_22,WX6176);
  and AND2_1849(WX5338,WX7540,WX5339);
  and AND2_1850(WX5341,WX5675,WX6176);
  and AND2_1851(WX5342,WX6247,WX5343);
  and AND2_1852(WX5347,WX5358,WX6175);
  and AND2_1853(WX5348,WX5354,WX5349);
  and AND2_1854(WX5351,CRC_OUT_5_21,WX6176);
  and AND2_1855(WX5352,WX7547,WX5353);
  and AND2_1856(WX5355,WX5677,WX6176);
  and AND2_1857(WX5356,WX6254,WX5357);
  and AND2_1858(WX5361,WX5372,WX6175);
  and AND2_1859(WX5362,WX5368,WX5363);
  and AND2_1860(WX5365,CRC_OUT_5_20,WX6176);
  and AND2_1861(WX5366,WX7554,WX5367);
  and AND2_1862(WX5369,WX5679,WX6176);
  and AND2_1863(WX5370,WX6261,WX5371);
  and AND2_1864(WX5375,WX5386,WX6175);
  and AND2_1865(WX5376,WX5382,WX5377);
  and AND2_1866(WX5379,CRC_OUT_5_19,WX6176);
  and AND2_1867(WX5380,WX7561,WX5381);
  and AND2_1868(WX5383,WX5681,WX6176);
  and AND2_1869(WX5384,WX6268,WX5385);
  and AND2_1870(WX5389,WX5400,WX6175);
  and AND2_1871(WX5390,WX5396,WX5391);
  and AND2_1872(WX5393,CRC_OUT_5_18,WX6176);
  and AND2_1873(WX5394,WX7568,WX5395);
  and AND2_1874(WX5397,WX5683,WX6176);
  and AND2_1875(WX5398,WX6275,WX5399);
  and AND2_1876(WX5403,WX5414,WX6175);
  and AND2_1877(WX5404,WX5410,WX5405);
  and AND2_1878(WX5407,CRC_OUT_5_17,WX6176);
  and AND2_1879(WX5408,WX7575,WX5409);
  and AND2_1880(WX5411,WX5685,WX6176);
  and AND2_1881(WX5412,WX6282,WX5413);
  and AND2_1882(WX5417,WX5428,WX6175);
  and AND2_1883(WX5418,WX5424,WX5419);
  and AND2_1884(WX5421,CRC_OUT_5_16,WX6176);
  and AND2_1885(WX5422,WX7582,WX5423);
  and AND2_1886(WX5425,WX5687,WX6176);
  and AND2_1887(WX5426,WX6289,WX5427);
  and AND2_1888(WX5431,WX5442,WX6175);
  and AND2_1889(WX5432,WX5438,WX5433);
  and AND2_1890(WX5435,CRC_OUT_5_15,WX6176);
  and AND2_1891(WX5436,WX7589,WX5437);
  and AND2_1892(WX5439,WX5689,WX6176);
  and AND2_1893(WX5440,WX6296,WX5441);
  and AND2_1894(WX5445,WX5456,WX6175);
  and AND2_1895(WX5446,WX5452,WX5447);
  and AND2_1896(WX5449,CRC_OUT_5_14,WX6176);
  and AND2_1897(WX5450,WX7596,WX5451);
  and AND2_1898(WX5453,WX5691,WX6176);
  and AND2_1899(WX5454,WX6303,WX5455);
  and AND2_1900(WX5459,WX5470,WX6175);
  and AND2_1901(WX5460,WX5466,WX5461);
  and AND2_1902(WX5463,CRC_OUT_5_13,WX6176);
  and AND2_1903(WX5464,WX7603,WX5465);
  and AND2_1904(WX5467,WX5693,WX6176);
  and AND2_1905(WX5468,WX6310,WX5469);
  and AND2_1906(WX5473,WX5484,WX6175);
  and AND2_1907(WX5474,WX5480,WX5475);
  and AND2_1908(WX5477,CRC_OUT_5_12,WX6176);
  and AND2_1909(WX5478,WX7610,WX5479);
  and AND2_1910(WX5481,WX5695,WX6176);
  and AND2_1911(WX5482,WX6317,WX5483);
  and AND2_1912(WX5487,WX5498,WX6175);
  and AND2_1913(WX5488,WX5494,WX5489);
  and AND2_1914(WX5491,CRC_OUT_5_11,WX6176);
  and AND2_1915(WX5492,WX7617,WX5493);
  and AND2_1916(WX5495,WX5697,WX6176);
  and AND2_1917(WX5496,WX6324,WX5497);
  and AND2_1918(WX5501,WX5512,WX6175);
  and AND2_1919(WX5502,WX5508,WX5503);
  and AND2_1920(WX5505,CRC_OUT_5_10,WX6176);
  and AND2_1921(WX5506,WX7624,WX5507);
  and AND2_1922(WX5509,WX5699,WX6176);
  and AND2_1923(WX5510,WX6331,WX5511);
  and AND2_1924(WX5515,WX5526,WX6175);
  and AND2_1925(WX5516,WX5522,WX5517);
  and AND2_1926(WX5519,CRC_OUT_5_9,WX6176);
  and AND2_1927(WX5520,WX7631,WX5521);
  and AND2_1928(WX5523,WX5701,WX6176);
  and AND2_1929(WX5524,WX6338,WX5525);
  and AND2_1930(WX5529,WX5540,WX6175);
  and AND2_1931(WX5530,WX5536,WX5531);
  and AND2_1932(WX5533,CRC_OUT_5_8,WX6176);
  and AND2_1933(WX5534,WX7638,WX5535);
  and AND2_1934(WX5537,WX5703,WX6176);
  and AND2_1935(WX5538,WX6345,WX5539);
  and AND2_1936(WX5543,WX5554,WX6175);
  and AND2_1937(WX5544,WX5550,WX5545);
  and AND2_1938(WX5547,CRC_OUT_5_7,WX6176);
  and AND2_1939(WX5548,WX7645,WX5549);
  and AND2_1940(WX5551,WX5705,WX6176);
  and AND2_1941(WX5552,WX6352,WX5553);
  and AND2_1942(WX5557,WX5568,WX6175);
  and AND2_1943(WX5558,WX5564,WX5559);
  and AND2_1944(WX5561,CRC_OUT_5_6,WX6176);
  and AND2_1945(WX5562,WX7652,WX5563);
  and AND2_1946(WX5565,WX5707,WX6176);
  and AND2_1947(WX5566,WX6359,WX5567);
  and AND2_1948(WX5571,WX5582,WX6175);
  and AND2_1949(WX5572,WX5578,WX5573);
  and AND2_1950(WX5575,CRC_OUT_5_5,WX6176);
  and AND2_1951(WX5576,WX7659,WX5577);
  and AND2_1952(WX5579,WX5709,WX6176);
  and AND2_1953(WX5580,WX6366,WX5581);
  and AND2_1954(WX5585,WX5596,WX6175);
  and AND2_1955(WX5586,WX5592,WX5587);
  and AND2_1956(WX5589,CRC_OUT_5_4,WX6176);
  and AND2_1957(WX5590,WX7666,WX5591);
  and AND2_1958(WX5593,WX5711,WX6176);
  and AND2_1959(WX5594,WX6373,WX5595);
  and AND2_1960(WX5599,WX5610,WX6175);
  and AND2_1961(WX5600,WX5606,WX5601);
  and AND2_1962(WX5603,CRC_OUT_5_3,WX6176);
  and AND2_1963(WX5604,WX7673,WX5605);
  and AND2_1964(WX5607,WX5713,WX6176);
  and AND2_1965(WX5608,WX6380,WX5609);
  and AND2_1966(WX5613,WX5624,WX6175);
  and AND2_1967(WX5614,WX5620,WX5615);
  and AND2_1968(WX5617,CRC_OUT_5_2,WX6176);
  and AND2_1969(WX5618,WX7680,WX5619);
  and AND2_1970(WX5621,WX5715,WX6176);
  and AND2_1971(WX5622,WX6387,WX5623);
  and AND2_1972(WX5627,WX5638,WX6175);
  and AND2_1973(WX5628,WX5634,WX5629);
  and AND2_1974(WX5631,CRC_OUT_5_1,WX6176);
  and AND2_1975(WX5632,WX7687,WX5633);
  and AND2_1976(WX5635,WX5717,WX6176);
  and AND2_1977(WX5636,WX6394,WX5637);
  and AND2_1978(WX5641,WX5652,WX6175);
  and AND2_1979(WX5642,WX5648,WX5643);
  and AND2_1980(WX5645,CRC_OUT_5_0,WX6176);
  and AND2_1981(WX5646,WX7694,WX5647);
  and AND2_1982(WX5649,WX5719,WX6176);
  and AND2_1983(WX5650,WX6401,WX5651);
  and AND2_1984(WX5656,WX5659,RESET);
  and AND2_1985(WX5658,WX5661,RESET);
  and AND2_1986(WX5660,WX5663,RESET);
  and AND2_1987(WX5662,WX5665,RESET);
  and AND2_1988(WX5664,WX5667,RESET);
  and AND2_1989(WX5666,WX5669,RESET);
  and AND2_1990(WX5668,WX5671,RESET);
  and AND2_1991(WX5670,WX5673,RESET);
  and AND2_1992(WX5672,WX5675,RESET);
  and AND2_1993(WX5674,WX5677,RESET);
  and AND2_1994(WX5676,WX5679,RESET);
  and AND2_1995(WX5678,WX5681,RESET);
  and AND2_1996(WX5680,WX5683,RESET);
  and AND2_1997(WX5682,WX5685,RESET);
  and AND2_1998(WX5684,WX5687,RESET);
  and AND2_1999(WX5686,WX5689,RESET);
  and AND2_2000(WX5688,WX5691,RESET);
  and AND2_2001(WX5690,WX5693,RESET);
  and AND2_2002(WX5692,WX5695,RESET);
  and AND2_2003(WX5694,WX5697,RESET);
  and AND2_2004(WX5696,WX5699,RESET);
  and AND2_2005(WX5698,WX5701,RESET);
  and AND2_2006(WX5700,WX5703,RESET);
  and AND2_2007(WX5702,WX5705,RESET);
  and AND2_2008(WX5704,WX5707,RESET);
  and AND2_2009(WX5706,WX5709,RESET);
  and AND2_2010(WX5708,WX5711,RESET);
  and AND2_2011(WX5710,WX5713,RESET);
  and AND2_2012(WX5712,WX5715,RESET);
  and AND2_2013(WX5714,WX5717,RESET);
  and AND2_2014(WX5716,WX5719,RESET);
  and AND2_2015(WX5718,WX5655,RESET);
  and AND2_2016(WX5816,WX5220,RESET);
  and AND2_2017(WX5818,WX5234,RESET);
  and AND2_2018(WX5820,WX5248,RESET);
  and AND2_2019(WX5822,WX5262,RESET);
  and AND2_2020(WX5824,WX5276,RESET);
  and AND2_2021(WX5826,WX5290,RESET);
  and AND2_2022(WX5828,WX5304,RESET);
  and AND2_2023(WX5830,WX5318,RESET);
  and AND2_2024(WX5832,WX5332,RESET);
  and AND2_2025(WX5834,WX5346,RESET);
  and AND2_2026(WX5836,WX5360,RESET);
  and AND2_2027(WX5838,WX5374,RESET);
  and AND2_2028(WX5840,WX5388,RESET);
  and AND2_2029(WX5842,WX5402,RESET);
  and AND2_2030(WX5844,WX5416,RESET);
  and AND2_2031(WX5846,WX5430,RESET);
  and AND2_2032(WX5848,WX5444,RESET);
  and AND2_2033(WX5850,WX5458,RESET);
  and AND2_2034(WX5852,WX5472,RESET);
  and AND2_2035(WX5854,WX5486,RESET);
  and AND2_2036(WX5856,WX5500,RESET);
  and AND2_2037(WX5858,WX5514,RESET);
  and AND2_2038(WX5860,WX5528,RESET);
  and AND2_2039(WX5862,WX5542,RESET);
  and AND2_2040(WX5864,WX5556,RESET);
  and AND2_2041(WX5866,WX5570,RESET);
  and AND2_2042(WX5868,WX5584,RESET);
  and AND2_2043(WX5870,WX5598,RESET);
  and AND2_2044(WX5872,WX5612,RESET);
  and AND2_2045(WX5874,WX5626,RESET);
  and AND2_2046(WX5876,WX5640,RESET);
  and AND2_2047(WX5878,WX5654,RESET);
  and AND2_2048(WX5880,WX5817,RESET);
  and AND2_2049(WX5882,WX5819,RESET);
  and AND2_2050(WX5884,WX5821,RESET);
  and AND2_2051(WX5886,WX5823,RESET);
  and AND2_2052(WX5888,WX5825,RESET);
  and AND2_2053(WX5890,WX5827,RESET);
  and AND2_2054(WX5892,WX5829,RESET);
  and AND2_2055(WX5894,WX5831,RESET);
  and AND2_2056(WX5896,WX5833,RESET);
  and AND2_2057(WX5898,WX5835,RESET);
  and AND2_2058(WX5900,WX5837,RESET);
  and AND2_2059(WX5902,WX5839,RESET);
  and AND2_2060(WX5904,WX5841,RESET);
  and AND2_2061(WX5906,WX5843,RESET);
  and AND2_2062(WX5908,WX5845,RESET);
  and AND2_2063(WX5910,WX5847,RESET);
  and AND2_2064(WX5912,WX5849,RESET);
  and AND2_2065(WX5914,WX5851,RESET);
  and AND2_2066(WX5916,WX5853,RESET);
  and AND2_2067(WX5918,WX5855,RESET);
  and AND2_2068(WX5920,WX5857,RESET);
  and AND2_2069(WX5922,WX5859,RESET);
  and AND2_2070(WX5924,WX5861,RESET);
  and AND2_2071(WX5926,WX5863,RESET);
  and AND2_2072(WX5928,WX5865,RESET);
  and AND2_2073(WX5930,WX5867,RESET);
  and AND2_2074(WX5932,WX5869,RESET);
  and AND2_2075(WX5934,WX5871,RESET);
  and AND2_2076(WX5936,WX5873,RESET);
  and AND2_2077(WX5938,WX5875,RESET);
  and AND2_2078(WX5940,WX5877,RESET);
  and AND2_2079(WX5942,WX5879,RESET);
  and AND2_2080(WX5944,WX5881,RESET);
  and AND2_2081(WX5946,WX5883,RESET);
  and AND2_2082(WX5948,WX5885,RESET);
  and AND2_2083(WX5950,WX5887,RESET);
  and AND2_2084(WX5952,WX5889,RESET);
  and AND2_2085(WX5954,WX5891,RESET);
  and AND2_2086(WX5956,WX5893,RESET);
  and AND2_2087(WX5958,WX5895,RESET);
  and AND2_2088(WX5960,WX5897,RESET);
  and AND2_2089(WX5962,WX5899,RESET);
  and AND2_2090(WX5964,WX5901,RESET);
  and AND2_2091(WX5966,WX5903,RESET);
  and AND2_2092(WX5968,WX5905,RESET);
  and AND2_2093(WX5970,WX5907,RESET);
  and AND2_2094(WX5972,WX5909,RESET);
  and AND2_2095(WX5974,WX5911,RESET);
  and AND2_2096(WX5976,WX5913,RESET);
  and AND2_2097(WX5978,WX5915,RESET);
  and AND2_2098(WX5980,WX5917,RESET);
  and AND2_2099(WX5982,WX5919,RESET);
  and AND2_2100(WX5984,WX5921,RESET);
  and AND2_2101(WX5986,WX5923,RESET);
  and AND2_2102(WX5988,WX5925,RESET);
  and AND2_2103(WX5990,WX5927,RESET);
  and AND2_2104(WX5992,WX5929,RESET);
  and AND2_2105(WX5994,WX5931,RESET);
  and AND2_2106(WX5996,WX5933,RESET);
  and AND2_2107(WX5998,WX5935,RESET);
  and AND2_2108(WX6000,WX5937,RESET);
  and AND2_2109(WX6002,WX5939,RESET);
  and AND2_2110(WX6004,WX5941,RESET);
  and AND2_2111(WX6006,WX5943,RESET);
  and AND2_2112(WX6008,WX5945,RESET);
  and AND2_2113(WX6010,WX5947,RESET);
  and AND2_2114(WX6012,WX5949,RESET);
  and AND2_2115(WX6014,WX5951,RESET);
  and AND2_2116(WX6016,WX5953,RESET);
  and AND2_2117(WX6018,WX5955,RESET);
  and AND2_2118(WX6020,WX5957,RESET);
  and AND2_2119(WX6022,WX5959,RESET);
  and AND2_2120(WX6024,WX5961,RESET);
  and AND2_2121(WX6026,WX5963,RESET);
  and AND2_2122(WX6028,WX5965,RESET);
  and AND2_2123(WX6030,WX5967,RESET);
  and AND2_2124(WX6032,WX5969,RESET);
  and AND2_2125(WX6034,WX5971,RESET);
  and AND2_2126(WX6036,WX5973,RESET);
  and AND2_2127(WX6038,WX5975,RESET);
  and AND2_2128(WX6040,WX5977,RESET);
  and AND2_2129(WX6042,WX5979,RESET);
  and AND2_2130(WX6044,WX5981,RESET);
  and AND2_2131(WX6046,WX5983,RESET);
  and AND2_2132(WX6048,WX5985,RESET);
  and AND2_2133(WX6050,WX5987,RESET);
  and AND2_2134(WX6052,WX5989,RESET);
  and AND2_2135(WX6054,WX5991,RESET);
  and AND2_2136(WX6056,WX5993,RESET);
  and AND2_2137(WX6058,WX5995,RESET);
  and AND2_2138(WX6060,WX5997,RESET);
  and AND2_2139(WX6062,WX5999,RESET);
  and AND2_2140(WX6064,WX6001,RESET);
  and AND2_2141(WX6066,WX6003,RESET);
  and AND2_2142(WX6068,WX6005,RESET);
  and AND2_2143(WX6070,WX6007,RESET);
  and AND2_2144(WX6179,WX6178,WX6177);
  and AND2_2145(WX6180,WX5752,WX6181);
  and AND2_2146(WX6186,WX6185,WX6177);
  and AND2_2147(WX6187,WX5753,WX6188);
  and AND2_2148(WX6193,WX6192,WX6177);
  and AND2_2149(WX6194,WX5754,WX6195);
  and AND2_2150(WX6200,WX6199,WX6177);
  and AND2_2151(WX6201,WX5755,WX6202);
  and AND2_2152(WX6207,WX6206,WX6177);
  and AND2_2153(WX6208,WX5756,WX6209);
  and AND2_2154(WX6214,WX6213,WX6177);
  and AND2_2155(WX6215,WX5757,WX6216);
  and AND2_2156(WX6221,WX6220,WX6177);
  and AND2_2157(WX6222,WX5758,WX6223);
  and AND2_2158(WX6228,WX6227,WX6177);
  and AND2_2159(WX6229,WX5759,WX6230);
  and AND2_2160(WX6235,WX6234,WX6177);
  and AND2_2161(WX6236,WX5760,WX6237);
  and AND2_2162(WX6242,WX6241,WX6177);
  and AND2_2163(WX6243,WX5761,WX6244);
  and AND2_2164(WX6249,WX6248,WX6177);
  and AND2_2165(WX6250,WX5762,WX6251);
  and AND2_2166(WX6256,WX6255,WX6177);
  and AND2_2167(WX6257,WX5763,WX6258);
  and AND2_2168(WX6263,WX6262,WX6177);
  and AND2_2169(WX6264,WX5764,WX6265);
  and AND2_2170(WX6270,WX6269,WX6177);
  and AND2_2171(WX6271,WX5765,WX6272);
  and AND2_2172(WX6277,WX6276,WX6177);
  and AND2_2173(WX6278,WX5766,WX6279);
  and AND2_2174(WX6284,WX6283,WX6177);
  and AND2_2175(WX6285,WX5767,WX6286);
  and AND2_2176(WX6291,WX6290,WX6177);
  and AND2_2177(WX6292,WX5768,WX6293);
  and AND2_2178(WX6298,WX6297,WX6177);
  and AND2_2179(WX6299,WX5769,WX6300);
  and AND2_2180(WX6305,WX6304,WX6177);
  and AND2_2181(WX6306,WX5770,WX6307);
  and AND2_2182(WX6312,WX6311,WX6177);
  and AND2_2183(WX6313,WX5771,WX6314);
  and AND2_2184(WX6319,WX6318,WX6177);
  and AND2_2185(WX6320,WX5772,WX6321);
  and AND2_2186(WX6326,WX6325,WX6177);
  and AND2_2187(WX6327,WX5773,WX6328);
  and AND2_2188(WX6333,WX6332,WX6177);
  and AND2_2189(WX6334,WX5774,WX6335);
  and AND2_2190(WX6340,WX6339,WX6177);
  and AND2_2191(WX6341,WX5775,WX6342);
  and AND2_2192(WX6347,WX6346,WX6177);
  and AND2_2193(WX6348,WX5776,WX6349);
  and AND2_2194(WX6354,WX6353,WX6177);
  and AND2_2195(WX6355,WX5777,WX6356);
  and AND2_2196(WX6361,WX6360,WX6177);
  and AND2_2197(WX6362,WX5778,WX6363);
  and AND2_2198(WX6368,WX6367,WX6177);
  and AND2_2199(WX6369,WX5779,WX6370);
  and AND2_2200(WX6375,WX6374,WX6177);
  and AND2_2201(WX6376,WX5780,WX6377);
  and AND2_2202(WX6382,WX6381,WX6177);
  and AND2_2203(WX6383,WX5781,WX6384);
  and AND2_2204(WX6389,WX6388,WX6177);
  and AND2_2205(WX6390,WX5782,WX6391);
  and AND2_2206(WX6396,WX6395,WX6177);
  and AND2_2207(WX6397,WX5783,WX6398);
  and AND2_2208(WX6436,WX6406,WX6435);
  and AND2_2209(WX6438,WX6434,WX6435);
  and AND2_2210(WX6440,WX6433,WX6435);
  and AND2_2211(WX6442,WX6432,WX6435);
  and AND2_2212(WX6444,WX6405,WX6435);
  and AND2_2213(WX6446,WX6431,WX6435);
  and AND2_2214(WX6448,WX6430,WX6435);
  and AND2_2215(WX6450,WX6429,WX6435);
  and AND2_2216(WX6452,WX6428,WX6435);
  and AND2_2217(WX6454,WX6427,WX6435);
  and AND2_2218(WX6456,WX6426,WX6435);
  and AND2_2219(WX6458,WX6404,WX6435);
  and AND2_2220(WX6460,WX6425,WX6435);
  and AND2_2221(WX6462,WX6424,WX6435);
  and AND2_2222(WX6464,WX6423,WX6435);
  and AND2_2223(WX6466,WX6422,WX6435);
  and AND2_2224(WX6468,WX6403,WX6435);
  and AND2_2225(WX6470,WX6421,WX6435);
  and AND2_2226(WX6472,WX6420,WX6435);
  and AND2_2227(WX6474,WX6419,WX6435);
  and AND2_2228(WX6476,WX6418,WX6435);
  and AND2_2229(WX6478,WX6417,WX6435);
  and AND2_2230(WX6480,WX6416,WX6435);
  and AND2_2231(WX6482,WX6415,WX6435);
  and AND2_2232(WX6484,WX6414,WX6435);
  and AND2_2233(WX6486,WX6413,WX6435);
  and AND2_2234(WX6488,WX6412,WX6435);
  and AND2_2235(WX6490,WX6411,WX6435);
  and AND2_2236(WX6492,WX6410,WX6435);
  and AND2_2237(WX6494,WX6409,WX6435);
  and AND2_2238(WX6496,WX6408,WX6435);
  and AND2_2239(WX6498,WX6407,WX6435);
  and AND2_2240(WX6500,WX6511,WX7468);
  and AND2_2241(WX6501,WX6507,WX6502);
  and AND2_2242(WX6504,CRC_OUT_4_31,WX7469);
  and AND2_2243(WX6505,WX8770,WX6506);
  and AND2_2244(WX6508,WX6950,WX7469);
  and AND2_2245(WX6509,WX7477,WX6510);
  and AND2_2246(WX6514,WX6525,WX7468);
  and AND2_2247(WX6515,WX6521,WX6516);
  and AND2_2248(WX6518,CRC_OUT_4_30,WX7469);
  and AND2_2249(WX6519,WX8777,WX6520);
  and AND2_2250(WX6522,WX6952,WX7469);
  and AND2_2251(WX6523,WX7484,WX6524);
  and AND2_2252(WX6528,WX6539,WX7468);
  and AND2_2253(WX6529,WX6535,WX6530);
  and AND2_2254(WX6532,CRC_OUT_4_29,WX7469);
  and AND2_2255(WX6533,WX8784,WX6534);
  and AND2_2256(WX6536,WX6954,WX7469);
  and AND2_2257(WX6537,WX7491,WX6538);
  and AND2_2258(WX6542,WX6553,WX7468);
  and AND2_2259(WX6543,WX6549,WX6544);
  and AND2_2260(WX6546,CRC_OUT_4_28,WX7469);
  and AND2_2261(WX6547,WX8791,WX6548);
  and AND2_2262(WX6550,WX6956,WX7469);
  and AND2_2263(WX6551,WX7498,WX6552);
  and AND2_2264(WX6556,WX6567,WX7468);
  and AND2_2265(WX6557,WX6563,WX6558);
  and AND2_2266(WX6560,CRC_OUT_4_27,WX7469);
  and AND2_2267(WX6561,WX8798,WX6562);
  and AND2_2268(WX6564,WX6958,WX7469);
  and AND2_2269(WX6565,WX7505,WX6566);
  and AND2_2270(WX6570,WX6581,WX7468);
  and AND2_2271(WX6571,WX6577,WX6572);
  and AND2_2272(WX6574,CRC_OUT_4_26,WX7469);
  and AND2_2273(WX6575,WX8805,WX6576);
  and AND2_2274(WX6578,WX6960,WX7469);
  and AND2_2275(WX6579,WX7512,WX6580);
  and AND2_2276(WX6584,WX6595,WX7468);
  and AND2_2277(WX6585,WX6591,WX6586);
  and AND2_2278(WX6588,CRC_OUT_4_25,WX7469);
  and AND2_2279(WX6589,WX8812,WX6590);
  and AND2_2280(WX6592,WX6962,WX7469);
  and AND2_2281(WX6593,WX7519,WX6594);
  and AND2_2282(WX6598,WX6609,WX7468);
  and AND2_2283(WX6599,WX6605,WX6600);
  and AND2_2284(WX6602,CRC_OUT_4_24,WX7469);
  and AND2_2285(WX6603,WX8819,WX6604);
  and AND2_2286(WX6606,WX6964,WX7469);
  and AND2_2287(WX6607,WX7526,WX6608);
  and AND2_2288(WX6612,WX6623,WX7468);
  and AND2_2289(WX6613,WX6619,WX6614);
  and AND2_2290(WX6616,CRC_OUT_4_23,WX7469);
  and AND2_2291(WX6617,WX8826,WX6618);
  and AND2_2292(WX6620,WX6966,WX7469);
  and AND2_2293(WX6621,WX7533,WX6622);
  and AND2_2294(WX6626,WX6637,WX7468);
  and AND2_2295(WX6627,WX6633,WX6628);
  and AND2_2296(WX6630,CRC_OUT_4_22,WX7469);
  and AND2_2297(WX6631,WX8833,WX6632);
  and AND2_2298(WX6634,WX6968,WX7469);
  and AND2_2299(WX6635,WX7540,WX6636);
  and AND2_2300(WX6640,WX6651,WX7468);
  and AND2_2301(WX6641,WX6647,WX6642);
  and AND2_2302(WX6644,CRC_OUT_4_21,WX7469);
  and AND2_2303(WX6645,WX8840,WX6646);
  and AND2_2304(WX6648,WX6970,WX7469);
  and AND2_2305(WX6649,WX7547,WX6650);
  and AND2_2306(WX6654,WX6665,WX7468);
  and AND2_2307(WX6655,WX6661,WX6656);
  and AND2_2308(WX6658,CRC_OUT_4_20,WX7469);
  and AND2_2309(WX6659,WX8847,WX6660);
  and AND2_2310(WX6662,WX6972,WX7469);
  and AND2_2311(WX6663,WX7554,WX6664);
  and AND2_2312(WX6668,WX6679,WX7468);
  and AND2_2313(WX6669,WX6675,WX6670);
  and AND2_2314(WX6672,CRC_OUT_4_19,WX7469);
  and AND2_2315(WX6673,WX8854,WX6674);
  and AND2_2316(WX6676,WX6974,WX7469);
  and AND2_2317(WX6677,WX7561,WX6678);
  and AND2_2318(WX6682,WX6693,WX7468);
  and AND2_2319(WX6683,WX6689,WX6684);
  and AND2_2320(WX6686,CRC_OUT_4_18,WX7469);
  and AND2_2321(WX6687,WX8861,WX6688);
  and AND2_2322(WX6690,WX6976,WX7469);
  and AND2_2323(WX6691,WX7568,WX6692);
  and AND2_2324(WX6696,WX6707,WX7468);
  and AND2_2325(WX6697,WX6703,WX6698);
  and AND2_2326(WX6700,CRC_OUT_4_17,WX7469);
  and AND2_2327(WX6701,WX8868,WX6702);
  and AND2_2328(WX6704,WX6978,WX7469);
  and AND2_2329(WX6705,WX7575,WX6706);
  and AND2_2330(WX6710,WX6721,WX7468);
  and AND2_2331(WX6711,WX6717,WX6712);
  and AND2_2332(WX6714,CRC_OUT_4_16,WX7469);
  and AND2_2333(WX6715,WX8875,WX6716);
  and AND2_2334(WX6718,WX6980,WX7469);
  and AND2_2335(WX6719,WX7582,WX6720);
  and AND2_2336(WX6724,WX6735,WX7468);
  and AND2_2337(WX6725,WX6731,WX6726);
  and AND2_2338(WX6728,CRC_OUT_4_15,WX7469);
  and AND2_2339(WX6729,WX8882,WX6730);
  and AND2_2340(WX6732,WX6982,WX7469);
  and AND2_2341(WX6733,WX7589,WX6734);
  and AND2_2342(WX6738,WX6749,WX7468);
  and AND2_2343(WX6739,WX6745,WX6740);
  and AND2_2344(WX6742,CRC_OUT_4_14,WX7469);
  and AND2_2345(WX6743,WX8889,WX6744);
  and AND2_2346(WX6746,WX6984,WX7469);
  and AND2_2347(WX6747,WX7596,WX6748);
  and AND2_2348(WX6752,WX6763,WX7468);
  and AND2_2349(WX6753,WX6759,WX6754);
  and AND2_2350(WX6756,CRC_OUT_4_13,WX7469);
  and AND2_2351(WX6757,WX8896,WX6758);
  and AND2_2352(WX6760,WX6986,WX7469);
  and AND2_2353(WX6761,WX7603,WX6762);
  and AND2_2354(WX6766,WX6777,WX7468);
  and AND2_2355(WX6767,WX6773,WX6768);
  and AND2_2356(WX6770,CRC_OUT_4_12,WX7469);
  and AND2_2357(WX6771,WX8903,WX6772);
  and AND2_2358(WX6774,WX6988,WX7469);
  and AND2_2359(WX6775,WX7610,WX6776);
  and AND2_2360(WX6780,WX6791,WX7468);
  and AND2_2361(WX6781,WX6787,WX6782);
  and AND2_2362(WX6784,CRC_OUT_4_11,WX7469);
  and AND2_2363(WX6785,WX8910,WX6786);
  and AND2_2364(WX6788,WX6990,WX7469);
  and AND2_2365(WX6789,WX7617,WX6790);
  and AND2_2366(WX6794,WX6805,WX7468);
  and AND2_2367(WX6795,WX6801,WX6796);
  and AND2_2368(WX6798,CRC_OUT_4_10,WX7469);
  and AND2_2369(WX6799,WX8917,WX6800);
  and AND2_2370(WX6802,WX6992,WX7469);
  and AND2_2371(WX6803,WX7624,WX6804);
  and AND2_2372(WX6808,WX6819,WX7468);
  and AND2_2373(WX6809,WX6815,WX6810);
  and AND2_2374(WX6812,CRC_OUT_4_9,WX7469);
  and AND2_2375(WX6813,WX8924,WX6814);
  and AND2_2376(WX6816,WX6994,WX7469);
  and AND2_2377(WX6817,WX7631,WX6818);
  and AND2_2378(WX6822,WX6833,WX7468);
  and AND2_2379(WX6823,WX6829,WX6824);
  and AND2_2380(WX6826,CRC_OUT_4_8,WX7469);
  and AND2_2381(WX6827,WX8931,WX6828);
  and AND2_2382(WX6830,WX6996,WX7469);
  and AND2_2383(WX6831,WX7638,WX6832);
  and AND2_2384(WX6836,WX6847,WX7468);
  and AND2_2385(WX6837,WX6843,WX6838);
  and AND2_2386(WX6840,CRC_OUT_4_7,WX7469);
  and AND2_2387(WX6841,WX8938,WX6842);
  and AND2_2388(WX6844,WX6998,WX7469);
  and AND2_2389(WX6845,WX7645,WX6846);
  and AND2_2390(WX6850,WX6861,WX7468);
  and AND2_2391(WX6851,WX6857,WX6852);
  and AND2_2392(WX6854,CRC_OUT_4_6,WX7469);
  and AND2_2393(WX6855,WX8945,WX6856);
  and AND2_2394(WX6858,WX7000,WX7469);
  and AND2_2395(WX6859,WX7652,WX6860);
  and AND2_2396(WX6864,WX6875,WX7468);
  and AND2_2397(WX6865,WX6871,WX6866);
  and AND2_2398(WX6868,CRC_OUT_4_5,WX7469);
  and AND2_2399(WX6869,WX8952,WX6870);
  and AND2_2400(WX6872,WX7002,WX7469);
  and AND2_2401(WX6873,WX7659,WX6874);
  and AND2_2402(WX6878,WX6889,WX7468);
  and AND2_2403(WX6879,WX6885,WX6880);
  and AND2_2404(WX6882,CRC_OUT_4_4,WX7469);
  and AND2_2405(WX6883,WX8959,WX6884);
  and AND2_2406(WX6886,WX7004,WX7469);
  and AND2_2407(WX6887,WX7666,WX6888);
  and AND2_2408(WX6892,WX6903,WX7468);
  and AND2_2409(WX6893,WX6899,WX6894);
  and AND2_2410(WX6896,CRC_OUT_4_3,WX7469);
  and AND2_2411(WX6897,WX8966,WX6898);
  and AND2_2412(WX6900,WX7006,WX7469);
  and AND2_2413(WX6901,WX7673,WX6902);
  and AND2_2414(WX6906,WX6917,WX7468);
  and AND2_2415(WX6907,WX6913,WX6908);
  and AND2_2416(WX6910,CRC_OUT_4_2,WX7469);
  and AND2_2417(WX6911,WX8973,WX6912);
  and AND2_2418(WX6914,WX7008,WX7469);
  and AND2_2419(WX6915,WX7680,WX6916);
  and AND2_2420(WX6920,WX6931,WX7468);
  and AND2_2421(WX6921,WX6927,WX6922);
  and AND2_2422(WX6924,CRC_OUT_4_1,WX7469);
  and AND2_2423(WX6925,WX8980,WX6926);
  and AND2_2424(WX6928,WX7010,WX7469);
  and AND2_2425(WX6929,WX7687,WX6930);
  and AND2_2426(WX6934,WX6945,WX7468);
  and AND2_2427(WX6935,WX6941,WX6936);
  and AND2_2428(WX6938,CRC_OUT_4_0,WX7469);
  and AND2_2429(WX6939,WX8987,WX6940);
  and AND2_2430(WX6942,WX7012,WX7469);
  and AND2_2431(WX6943,WX7694,WX6944);
  and AND2_2432(WX6949,WX6952,RESET);
  and AND2_2433(WX6951,WX6954,RESET);
  and AND2_2434(WX6953,WX6956,RESET);
  and AND2_2435(WX6955,WX6958,RESET);
  and AND2_2436(WX6957,WX6960,RESET);
  and AND2_2437(WX6959,WX6962,RESET);
  and AND2_2438(WX6961,WX6964,RESET);
  and AND2_2439(WX6963,WX6966,RESET);
  and AND2_2440(WX6965,WX6968,RESET);
  and AND2_2441(WX6967,WX6970,RESET);
  and AND2_2442(WX6969,WX6972,RESET);
  and AND2_2443(WX6971,WX6974,RESET);
  and AND2_2444(WX6973,WX6976,RESET);
  and AND2_2445(WX6975,WX6978,RESET);
  and AND2_2446(WX6977,WX6980,RESET);
  and AND2_2447(WX6979,WX6982,RESET);
  and AND2_2448(WX6981,WX6984,RESET);
  and AND2_2449(WX6983,WX6986,RESET);
  and AND2_2450(WX6985,WX6988,RESET);
  and AND2_2451(WX6987,WX6990,RESET);
  and AND2_2452(WX6989,WX6992,RESET);
  and AND2_2453(WX6991,WX6994,RESET);
  and AND2_2454(WX6993,WX6996,RESET);
  and AND2_2455(WX6995,WX6998,RESET);
  and AND2_2456(WX6997,WX7000,RESET);
  and AND2_2457(WX6999,WX7002,RESET);
  and AND2_2458(WX7001,WX7004,RESET);
  and AND2_2459(WX7003,WX7006,RESET);
  and AND2_2460(WX7005,WX7008,RESET);
  and AND2_2461(WX7007,WX7010,RESET);
  and AND2_2462(WX7009,WX7012,RESET);
  and AND2_2463(WX7011,WX6948,RESET);
  and AND2_2464(WX7109,WX6513,RESET);
  and AND2_2465(WX7111,WX6527,RESET);
  and AND2_2466(WX7113,WX6541,RESET);
  and AND2_2467(WX7115,WX6555,RESET);
  and AND2_2468(WX7117,WX6569,RESET);
  and AND2_2469(WX7119,WX6583,RESET);
  and AND2_2470(WX7121,WX6597,RESET);
  and AND2_2471(WX7123,WX6611,RESET);
  and AND2_2472(WX7125,WX6625,RESET);
  and AND2_2473(WX7127,WX6639,RESET);
  and AND2_2474(WX7129,WX6653,RESET);
  and AND2_2475(WX7131,WX6667,RESET);
  and AND2_2476(WX7133,WX6681,RESET);
  and AND2_2477(WX7135,WX6695,RESET);
  and AND2_2478(WX7137,WX6709,RESET);
  and AND2_2479(WX7139,WX6723,RESET);
  and AND2_2480(WX7141,WX6737,RESET);
  and AND2_2481(WX7143,WX6751,RESET);
  and AND2_2482(WX7145,WX6765,RESET);
  and AND2_2483(WX7147,WX6779,RESET);
  and AND2_2484(WX7149,WX6793,RESET);
  and AND2_2485(WX7151,WX6807,RESET);
  and AND2_2486(WX7153,WX6821,RESET);
  and AND2_2487(WX7155,WX6835,RESET);
  and AND2_2488(WX7157,WX6849,RESET);
  and AND2_2489(WX7159,WX6863,RESET);
  and AND2_2490(WX7161,WX6877,RESET);
  and AND2_2491(WX7163,WX6891,RESET);
  and AND2_2492(WX7165,WX6905,RESET);
  and AND2_2493(WX7167,WX6919,RESET);
  and AND2_2494(WX7169,WX6933,RESET);
  and AND2_2495(WX7171,WX6947,RESET);
  and AND2_2496(WX7173,WX7110,RESET);
  and AND2_2497(WX7175,WX7112,RESET);
  and AND2_2498(WX7177,WX7114,RESET);
  and AND2_2499(WX7179,WX7116,RESET);
  and AND2_2500(WX7181,WX7118,RESET);
  and AND2_2501(WX7183,WX7120,RESET);
  and AND2_2502(WX7185,WX7122,RESET);
  and AND2_2503(WX7187,WX7124,RESET);
  and AND2_2504(WX7189,WX7126,RESET);
  and AND2_2505(WX7191,WX7128,RESET);
  and AND2_2506(WX7193,WX7130,RESET);
  and AND2_2507(WX7195,WX7132,RESET);
  and AND2_2508(WX7197,WX7134,RESET);
  and AND2_2509(WX7199,WX7136,RESET);
  and AND2_2510(WX7201,WX7138,RESET);
  and AND2_2511(WX7203,WX7140,RESET);
  and AND2_2512(WX7205,WX7142,RESET);
  and AND2_2513(WX7207,WX7144,RESET);
  and AND2_2514(WX7209,WX7146,RESET);
  and AND2_2515(WX7211,WX7148,RESET);
  and AND2_2516(WX7213,WX7150,RESET);
  and AND2_2517(WX7215,WX7152,RESET);
  and AND2_2518(WX7217,WX7154,RESET);
  and AND2_2519(WX7219,WX7156,RESET);
  and AND2_2520(WX7221,WX7158,RESET);
  and AND2_2521(WX7223,WX7160,RESET);
  and AND2_2522(WX7225,WX7162,RESET);
  and AND2_2523(WX7227,WX7164,RESET);
  and AND2_2524(WX7229,WX7166,RESET);
  and AND2_2525(WX7231,WX7168,RESET);
  and AND2_2526(WX7233,WX7170,RESET);
  and AND2_2527(WX7235,WX7172,RESET);
  and AND2_2528(WX7237,WX7174,RESET);
  and AND2_2529(WX7239,WX7176,RESET);
  and AND2_2530(WX7241,WX7178,RESET);
  and AND2_2531(WX7243,WX7180,RESET);
  and AND2_2532(WX7245,WX7182,RESET);
  and AND2_2533(WX7247,WX7184,RESET);
  and AND2_2534(WX7249,WX7186,RESET);
  and AND2_2535(WX7251,WX7188,RESET);
  and AND2_2536(WX7253,WX7190,RESET);
  and AND2_2537(WX7255,WX7192,RESET);
  and AND2_2538(WX7257,WX7194,RESET);
  and AND2_2539(WX7259,WX7196,RESET);
  and AND2_2540(WX7261,WX7198,RESET);
  and AND2_2541(WX7263,WX7200,RESET);
  and AND2_2542(WX7265,WX7202,RESET);
  and AND2_2543(WX7267,WX7204,RESET);
  and AND2_2544(WX7269,WX7206,RESET);
  and AND2_2545(WX7271,WX7208,RESET);
  and AND2_2546(WX7273,WX7210,RESET);
  and AND2_2547(WX7275,WX7212,RESET);
  and AND2_2548(WX7277,WX7214,RESET);
  and AND2_2549(WX7279,WX7216,RESET);
  and AND2_2550(WX7281,WX7218,RESET);
  and AND2_2551(WX7283,WX7220,RESET);
  and AND2_2552(WX7285,WX7222,RESET);
  and AND2_2553(WX7287,WX7224,RESET);
  and AND2_2554(WX7289,WX7226,RESET);
  and AND2_2555(WX7291,WX7228,RESET);
  and AND2_2556(WX7293,WX7230,RESET);
  and AND2_2557(WX7295,WX7232,RESET);
  and AND2_2558(WX7297,WX7234,RESET);
  and AND2_2559(WX7299,WX7236,RESET);
  and AND2_2560(WX7301,WX7238,RESET);
  and AND2_2561(WX7303,WX7240,RESET);
  and AND2_2562(WX7305,WX7242,RESET);
  and AND2_2563(WX7307,WX7244,RESET);
  and AND2_2564(WX7309,WX7246,RESET);
  and AND2_2565(WX7311,WX7248,RESET);
  and AND2_2566(WX7313,WX7250,RESET);
  and AND2_2567(WX7315,WX7252,RESET);
  and AND2_2568(WX7317,WX7254,RESET);
  and AND2_2569(WX7319,WX7256,RESET);
  and AND2_2570(WX7321,WX7258,RESET);
  and AND2_2571(WX7323,WX7260,RESET);
  and AND2_2572(WX7325,WX7262,RESET);
  and AND2_2573(WX7327,WX7264,RESET);
  and AND2_2574(WX7329,WX7266,RESET);
  and AND2_2575(WX7331,WX7268,RESET);
  and AND2_2576(WX7333,WX7270,RESET);
  and AND2_2577(WX7335,WX7272,RESET);
  and AND2_2578(WX7337,WX7274,RESET);
  and AND2_2579(WX7339,WX7276,RESET);
  and AND2_2580(WX7341,WX7278,RESET);
  and AND2_2581(WX7343,WX7280,RESET);
  and AND2_2582(WX7345,WX7282,RESET);
  and AND2_2583(WX7347,WX7284,RESET);
  and AND2_2584(WX7349,WX7286,RESET);
  and AND2_2585(WX7351,WX7288,RESET);
  and AND2_2586(WX7353,WX7290,RESET);
  and AND2_2587(WX7355,WX7292,RESET);
  and AND2_2588(WX7357,WX7294,RESET);
  and AND2_2589(WX7359,WX7296,RESET);
  and AND2_2590(WX7361,WX7298,RESET);
  and AND2_2591(WX7363,WX7300,RESET);
  and AND2_2592(WX7472,WX7471,WX7470);
  and AND2_2593(WX7473,WX7045,WX7474);
  and AND2_2594(WX7479,WX7478,WX7470);
  and AND2_2595(WX7480,WX7046,WX7481);
  and AND2_2596(WX7486,WX7485,WX7470);
  and AND2_2597(WX7487,WX7047,WX7488);
  and AND2_2598(WX7493,WX7492,WX7470);
  and AND2_2599(WX7494,WX7048,WX7495);
  and AND2_2600(WX7500,WX7499,WX7470);
  and AND2_2601(WX7501,WX7049,WX7502);
  and AND2_2602(WX7507,WX7506,WX7470);
  and AND2_2603(WX7508,WX7050,WX7509);
  and AND2_2604(WX7514,WX7513,WX7470);
  and AND2_2605(WX7515,WX7051,WX7516);
  and AND2_2606(WX7521,WX7520,WX7470);
  and AND2_2607(WX7522,WX7052,WX7523);
  and AND2_2608(WX7528,WX7527,WX7470);
  and AND2_2609(WX7529,WX7053,WX7530);
  and AND2_2610(WX7535,WX7534,WX7470);
  and AND2_2611(WX7536,WX7054,WX7537);
  and AND2_2612(WX7542,WX7541,WX7470);
  and AND2_2613(WX7543,WX7055,WX7544);
  and AND2_2614(WX7549,WX7548,WX7470);
  and AND2_2615(WX7550,WX7056,WX7551);
  and AND2_2616(WX7556,WX7555,WX7470);
  and AND2_2617(WX7557,WX7057,WX7558);
  and AND2_2618(WX7563,WX7562,WX7470);
  and AND2_2619(WX7564,WX7058,WX7565);
  and AND2_2620(WX7570,WX7569,WX7470);
  and AND2_2621(WX7571,WX7059,WX7572);
  and AND2_2622(WX7577,WX7576,WX7470);
  and AND2_2623(WX7578,WX7060,WX7579);
  and AND2_2624(WX7584,WX7583,WX7470);
  and AND2_2625(WX7585,WX7061,WX7586);
  and AND2_2626(WX7591,WX7590,WX7470);
  and AND2_2627(WX7592,WX7062,WX7593);
  and AND2_2628(WX7598,WX7597,WX7470);
  and AND2_2629(WX7599,WX7063,WX7600);
  and AND2_2630(WX7605,WX7604,WX7470);
  and AND2_2631(WX7606,WX7064,WX7607);
  and AND2_2632(WX7612,WX7611,WX7470);
  and AND2_2633(WX7613,WX7065,WX7614);
  and AND2_2634(WX7619,WX7618,WX7470);
  and AND2_2635(WX7620,WX7066,WX7621);
  and AND2_2636(WX7626,WX7625,WX7470);
  and AND2_2637(WX7627,WX7067,WX7628);
  and AND2_2638(WX7633,WX7632,WX7470);
  and AND2_2639(WX7634,WX7068,WX7635);
  and AND2_2640(WX7640,WX7639,WX7470);
  and AND2_2641(WX7641,WX7069,WX7642);
  and AND2_2642(WX7647,WX7646,WX7470);
  and AND2_2643(WX7648,WX7070,WX7649);
  and AND2_2644(WX7654,WX7653,WX7470);
  and AND2_2645(WX7655,WX7071,WX7656);
  and AND2_2646(WX7661,WX7660,WX7470);
  and AND2_2647(WX7662,WX7072,WX7663);
  and AND2_2648(WX7668,WX7667,WX7470);
  and AND2_2649(WX7669,WX7073,WX7670);
  and AND2_2650(WX7675,WX7674,WX7470);
  and AND2_2651(WX7676,WX7074,WX7677);
  and AND2_2652(WX7682,WX7681,WX7470);
  and AND2_2653(WX7683,WX7075,WX7684);
  and AND2_2654(WX7689,WX7688,WX7470);
  and AND2_2655(WX7690,WX7076,WX7691);
  and AND2_2656(WX7729,WX7699,WX7728);
  and AND2_2657(WX7731,WX7727,WX7728);
  and AND2_2658(WX7733,WX7726,WX7728);
  and AND2_2659(WX7735,WX7725,WX7728);
  and AND2_2660(WX7737,WX7698,WX7728);
  and AND2_2661(WX7739,WX7724,WX7728);
  and AND2_2662(WX7741,WX7723,WX7728);
  and AND2_2663(WX7743,WX7722,WX7728);
  and AND2_2664(WX7745,WX7721,WX7728);
  and AND2_2665(WX7747,WX7720,WX7728);
  and AND2_2666(WX7749,WX7719,WX7728);
  and AND2_2667(WX7751,WX7697,WX7728);
  and AND2_2668(WX7753,WX7718,WX7728);
  and AND2_2669(WX7755,WX7717,WX7728);
  and AND2_2670(WX7757,WX7716,WX7728);
  and AND2_2671(WX7759,WX7715,WX7728);
  and AND2_2672(WX7761,WX7696,WX7728);
  and AND2_2673(WX7763,WX7714,WX7728);
  and AND2_2674(WX7765,WX7713,WX7728);
  and AND2_2675(WX7767,WX7712,WX7728);
  and AND2_2676(WX7769,WX7711,WX7728);
  and AND2_2677(WX7771,WX7710,WX7728);
  and AND2_2678(WX7773,WX7709,WX7728);
  and AND2_2679(WX7775,WX7708,WX7728);
  and AND2_2680(WX7777,WX7707,WX7728);
  and AND2_2681(WX7779,WX7706,WX7728);
  and AND2_2682(WX7781,WX7705,WX7728);
  and AND2_2683(WX7783,WX7704,WX7728);
  and AND2_2684(WX7785,WX7703,WX7728);
  and AND2_2685(WX7787,WX7702,WX7728);
  and AND2_2686(WX7789,WX7701,WX7728);
  and AND2_2687(WX7791,WX7700,WX7728);
  and AND2_2688(WX7793,WX7804,WX8761);
  and AND2_2689(WX7794,WX7800,WX7795);
  and AND2_2690(WX7797,CRC_OUT_3_31,WX8762);
  and AND2_2691(WX7798,WX10063,WX7799);
  and AND2_2692(WX7801,WX8243,WX8762);
  and AND2_2693(WX7802,WX8770,WX7803);
  and AND2_2694(WX7807,WX7818,WX8761);
  and AND2_2695(WX7808,WX7814,WX7809);
  and AND2_2696(WX7811,CRC_OUT_3_30,WX8762);
  and AND2_2697(WX7812,WX10070,WX7813);
  and AND2_2698(WX7815,WX8245,WX8762);
  and AND2_2699(WX7816,WX8777,WX7817);
  and AND2_2700(WX7821,WX7832,WX8761);
  and AND2_2701(WX7822,WX7828,WX7823);
  and AND2_2702(WX7825,CRC_OUT_3_29,WX8762);
  and AND2_2703(WX7826,WX10077,WX7827);
  and AND2_2704(WX7829,WX8247,WX8762);
  and AND2_2705(WX7830,WX8784,WX7831);
  and AND2_2706(WX7835,WX7846,WX8761);
  and AND2_2707(WX7836,WX7842,WX7837);
  and AND2_2708(WX7839,CRC_OUT_3_28,WX8762);
  and AND2_2709(WX7840,WX10084,WX7841);
  and AND2_2710(WX7843,WX8249,WX8762);
  and AND2_2711(WX7844,WX8791,WX7845);
  and AND2_2712(WX7849,WX7860,WX8761);
  and AND2_2713(WX7850,WX7856,WX7851);
  and AND2_2714(WX7853,CRC_OUT_3_27,WX8762);
  and AND2_2715(WX7854,WX10091,WX7855);
  and AND2_2716(WX7857,WX8251,WX8762);
  and AND2_2717(WX7858,WX8798,WX7859);
  and AND2_2718(WX7863,WX7874,WX8761);
  and AND2_2719(WX7864,WX7870,WX7865);
  and AND2_2720(WX7867,CRC_OUT_3_26,WX8762);
  and AND2_2721(WX7868,WX10098,WX7869);
  and AND2_2722(WX7871,WX8253,WX8762);
  and AND2_2723(WX7872,WX8805,WX7873);
  and AND2_2724(WX7877,WX7888,WX8761);
  and AND2_2725(WX7878,WX7884,WX7879);
  and AND2_2726(WX7881,CRC_OUT_3_25,WX8762);
  and AND2_2727(WX7882,WX10105,WX7883);
  and AND2_2728(WX7885,WX8255,WX8762);
  and AND2_2729(WX7886,WX8812,WX7887);
  and AND2_2730(WX7891,WX7902,WX8761);
  and AND2_2731(WX7892,WX7898,WX7893);
  and AND2_2732(WX7895,CRC_OUT_3_24,WX8762);
  and AND2_2733(WX7896,WX10112,WX7897);
  and AND2_2734(WX7899,WX8257,WX8762);
  and AND2_2735(WX7900,WX8819,WX7901);
  and AND2_2736(WX7905,WX7916,WX8761);
  and AND2_2737(WX7906,WX7912,WX7907);
  and AND2_2738(WX7909,CRC_OUT_3_23,WX8762);
  and AND2_2739(WX7910,WX10119,WX7911);
  and AND2_2740(WX7913,WX8259,WX8762);
  and AND2_2741(WX7914,WX8826,WX7915);
  and AND2_2742(WX7919,WX7930,WX8761);
  and AND2_2743(WX7920,WX7926,WX7921);
  and AND2_2744(WX7923,CRC_OUT_3_22,WX8762);
  and AND2_2745(WX7924,WX10126,WX7925);
  and AND2_2746(WX7927,WX8261,WX8762);
  and AND2_2747(WX7928,WX8833,WX7929);
  and AND2_2748(WX7933,WX7944,WX8761);
  and AND2_2749(WX7934,WX7940,WX7935);
  and AND2_2750(WX7937,CRC_OUT_3_21,WX8762);
  and AND2_2751(WX7938,WX10133,WX7939);
  and AND2_2752(WX7941,WX8263,WX8762);
  and AND2_2753(WX7942,WX8840,WX7943);
  and AND2_2754(WX7947,WX7958,WX8761);
  and AND2_2755(WX7948,WX7954,WX7949);
  and AND2_2756(WX7951,CRC_OUT_3_20,WX8762);
  and AND2_2757(WX7952,WX10140,WX7953);
  and AND2_2758(WX7955,WX8265,WX8762);
  and AND2_2759(WX7956,WX8847,WX7957);
  and AND2_2760(WX7961,WX7972,WX8761);
  and AND2_2761(WX7962,WX7968,WX7963);
  and AND2_2762(WX7965,CRC_OUT_3_19,WX8762);
  and AND2_2763(WX7966,WX10147,WX7967);
  and AND2_2764(WX7969,WX8267,WX8762);
  and AND2_2765(WX7970,WX8854,WX7971);
  and AND2_2766(WX7975,WX7986,WX8761);
  and AND2_2767(WX7976,WX7982,WX7977);
  and AND2_2768(WX7979,CRC_OUT_3_18,WX8762);
  and AND2_2769(WX7980,WX10154,WX7981);
  and AND2_2770(WX7983,WX8269,WX8762);
  and AND2_2771(WX7984,WX8861,WX7985);
  and AND2_2772(WX7989,WX8000,WX8761);
  and AND2_2773(WX7990,WX7996,WX7991);
  and AND2_2774(WX7993,CRC_OUT_3_17,WX8762);
  and AND2_2775(WX7994,WX10161,WX7995);
  and AND2_2776(WX7997,WX8271,WX8762);
  and AND2_2777(WX7998,WX8868,WX7999);
  and AND2_2778(WX8003,WX8014,WX8761);
  and AND2_2779(WX8004,WX8010,WX8005);
  and AND2_2780(WX8007,CRC_OUT_3_16,WX8762);
  and AND2_2781(WX8008,WX10168,WX8009);
  and AND2_2782(WX8011,WX8273,WX8762);
  and AND2_2783(WX8012,WX8875,WX8013);
  and AND2_2784(WX8017,WX8028,WX8761);
  and AND2_2785(WX8018,WX8024,WX8019);
  and AND2_2786(WX8021,CRC_OUT_3_15,WX8762);
  and AND2_2787(WX8022,WX10175,WX8023);
  and AND2_2788(WX8025,WX8275,WX8762);
  and AND2_2789(WX8026,WX8882,WX8027);
  and AND2_2790(WX8031,WX8042,WX8761);
  and AND2_2791(WX8032,WX8038,WX8033);
  and AND2_2792(WX8035,CRC_OUT_3_14,WX8762);
  and AND2_2793(WX8036,WX10182,WX8037);
  and AND2_2794(WX8039,WX8277,WX8762);
  and AND2_2795(WX8040,WX8889,WX8041);
  and AND2_2796(WX8045,WX8056,WX8761);
  and AND2_2797(WX8046,WX8052,WX8047);
  and AND2_2798(WX8049,CRC_OUT_3_13,WX8762);
  and AND2_2799(WX8050,WX10189,WX8051);
  and AND2_2800(WX8053,WX8279,WX8762);
  and AND2_2801(WX8054,WX8896,WX8055);
  and AND2_2802(WX8059,WX8070,WX8761);
  and AND2_2803(WX8060,WX8066,WX8061);
  and AND2_2804(WX8063,CRC_OUT_3_12,WX8762);
  and AND2_2805(WX8064,WX10196,WX8065);
  and AND2_2806(WX8067,WX8281,WX8762);
  and AND2_2807(WX8068,WX8903,WX8069);
  and AND2_2808(WX8073,WX8084,WX8761);
  and AND2_2809(WX8074,WX8080,WX8075);
  and AND2_2810(WX8077,CRC_OUT_3_11,WX8762);
  and AND2_2811(WX8078,WX10203,WX8079);
  and AND2_2812(WX8081,WX8283,WX8762);
  and AND2_2813(WX8082,WX8910,WX8083);
  and AND2_2814(WX8087,WX8098,WX8761);
  and AND2_2815(WX8088,WX8094,WX8089);
  and AND2_2816(WX8091,CRC_OUT_3_10,WX8762);
  and AND2_2817(WX8092,WX10210,WX8093);
  and AND2_2818(WX8095,WX8285,WX8762);
  and AND2_2819(WX8096,WX8917,WX8097);
  and AND2_2820(WX8101,WX8112,WX8761);
  and AND2_2821(WX8102,WX8108,WX8103);
  and AND2_2822(WX8105,CRC_OUT_3_9,WX8762);
  and AND2_2823(WX8106,WX10217,WX8107);
  and AND2_2824(WX8109,WX8287,WX8762);
  and AND2_2825(WX8110,WX8924,WX8111);
  and AND2_2826(WX8115,WX8126,WX8761);
  and AND2_2827(WX8116,WX8122,WX8117);
  and AND2_2828(WX8119,CRC_OUT_3_8,WX8762);
  and AND2_2829(WX8120,WX10224,WX8121);
  and AND2_2830(WX8123,WX8289,WX8762);
  and AND2_2831(WX8124,WX8931,WX8125);
  and AND2_2832(WX8129,WX8140,WX8761);
  and AND2_2833(WX8130,WX8136,WX8131);
  and AND2_2834(WX8133,CRC_OUT_3_7,WX8762);
  and AND2_2835(WX8134,WX10231,WX8135);
  and AND2_2836(WX8137,WX8291,WX8762);
  and AND2_2837(WX8138,WX8938,WX8139);
  and AND2_2838(WX8143,WX8154,WX8761);
  and AND2_2839(WX8144,WX8150,WX8145);
  and AND2_2840(WX8147,CRC_OUT_3_6,WX8762);
  and AND2_2841(WX8148,WX10238,WX8149);
  and AND2_2842(WX8151,WX8293,WX8762);
  and AND2_2843(WX8152,WX8945,WX8153);
  and AND2_2844(WX8157,WX8168,WX8761);
  and AND2_2845(WX8158,WX8164,WX8159);
  and AND2_2846(WX8161,CRC_OUT_3_5,WX8762);
  and AND2_2847(WX8162,WX10245,WX8163);
  and AND2_2848(WX8165,WX8295,WX8762);
  and AND2_2849(WX8166,WX8952,WX8167);
  and AND2_2850(WX8171,WX8182,WX8761);
  and AND2_2851(WX8172,WX8178,WX8173);
  and AND2_2852(WX8175,CRC_OUT_3_4,WX8762);
  and AND2_2853(WX8176,WX10252,WX8177);
  and AND2_2854(WX8179,WX8297,WX8762);
  and AND2_2855(WX8180,WX8959,WX8181);
  and AND2_2856(WX8185,WX8196,WX8761);
  and AND2_2857(WX8186,WX8192,WX8187);
  and AND2_2858(WX8189,CRC_OUT_3_3,WX8762);
  and AND2_2859(WX8190,WX10259,WX8191);
  and AND2_2860(WX8193,WX8299,WX8762);
  and AND2_2861(WX8194,WX8966,WX8195);
  and AND2_2862(WX8199,WX8210,WX8761);
  and AND2_2863(WX8200,WX8206,WX8201);
  and AND2_2864(WX8203,CRC_OUT_3_2,WX8762);
  and AND2_2865(WX8204,WX10266,WX8205);
  and AND2_2866(WX8207,WX8301,WX8762);
  and AND2_2867(WX8208,WX8973,WX8209);
  and AND2_2868(WX8213,WX8224,WX8761);
  and AND2_2869(WX8214,WX8220,WX8215);
  and AND2_2870(WX8217,CRC_OUT_3_1,WX8762);
  and AND2_2871(WX8218,WX10273,WX8219);
  and AND2_2872(WX8221,WX8303,WX8762);
  and AND2_2873(WX8222,WX8980,WX8223);
  and AND2_2874(WX8227,WX8238,WX8761);
  and AND2_2875(WX8228,WX8234,WX8229);
  and AND2_2876(WX8231,CRC_OUT_3_0,WX8762);
  and AND2_2877(WX8232,WX10280,WX8233);
  and AND2_2878(WX8235,WX8305,WX8762);
  and AND2_2879(WX8236,WX8987,WX8237);
  and AND2_2880(WX8242,WX8245,RESET);
  and AND2_2881(WX8244,WX8247,RESET);
  and AND2_2882(WX8246,WX8249,RESET);
  and AND2_2883(WX8248,WX8251,RESET);
  and AND2_2884(WX8250,WX8253,RESET);
  and AND2_2885(WX8252,WX8255,RESET);
  and AND2_2886(WX8254,WX8257,RESET);
  and AND2_2887(WX8256,WX8259,RESET);
  and AND2_2888(WX8258,WX8261,RESET);
  and AND2_2889(WX8260,WX8263,RESET);
  and AND2_2890(WX8262,WX8265,RESET);
  and AND2_2891(WX8264,WX8267,RESET);
  and AND2_2892(WX8266,WX8269,RESET);
  and AND2_2893(WX8268,WX8271,RESET);
  and AND2_2894(WX8270,WX8273,RESET);
  and AND2_2895(WX8272,WX8275,RESET);
  and AND2_2896(WX8274,WX8277,RESET);
  and AND2_2897(WX8276,WX8279,RESET);
  and AND2_2898(WX8278,WX8281,RESET);
  and AND2_2899(WX8280,WX8283,RESET);
  and AND2_2900(WX8282,WX8285,RESET);
  and AND2_2901(WX8284,WX8287,RESET);
  and AND2_2902(WX8286,WX8289,RESET);
  and AND2_2903(WX8288,WX8291,RESET);
  and AND2_2904(WX8290,WX8293,RESET);
  and AND2_2905(WX8292,WX8295,RESET);
  and AND2_2906(WX8294,WX8297,RESET);
  and AND2_2907(WX8296,WX8299,RESET);
  and AND2_2908(WX8298,WX8301,RESET);
  and AND2_2909(WX8300,WX8303,RESET);
  and AND2_2910(WX8302,WX8305,RESET);
  and AND2_2911(WX8304,WX8241,RESET);
  and AND2_2912(WX8402,WX7806,RESET);
  and AND2_2913(WX8404,WX7820,RESET);
  and AND2_2914(WX8406,WX7834,RESET);
  and AND2_2915(WX8408,WX7848,RESET);
  and AND2_2916(WX8410,WX7862,RESET);
  and AND2_2917(WX8412,WX7876,RESET);
  and AND2_2918(WX8414,WX7890,RESET);
  and AND2_2919(WX8416,WX7904,RESET);
  and AND2_2920(WX8418,WX7918,RESET);
  and AND2_2921(WX8420,WX7932,RESET);
  and AND2_2922(WX8422,WX7946,RESET);
  and AND2_2923(WX8424,WX7960,RESET);
  and AND2_2924(WX8426,WX7974,RESET);
  and AND2_2925(WX8428,WX7988,RESET);
  and AND2_2926(WX8430,WX8002,RESET);
  and AND2_2927(WX8432,WX8016,RESET);
  and AND2_2928(WX8434,WX8030,RESET);
  and AND2_2929(WX8436,WX8044,RESET);
  and AND2_2930(WX8438,WX8058,RESET);
  and AND2_2931(WX8440,WX8072,RESET);
  and AND2_2932(WX8442,WX8086,RESET);
  and AND2_2933(WX8444,WX8100,RESET);
  and AND2_2934(WX8446,WX8114,RESET);
  and AND2_2935(WX8448,WX8128,RESET);
  and AND2_2936(WX8450,WX8142,RESET);
  and AND2_2937(WX8452,WX8156,RESET);
  and AND2_2938(WX8454,WX8170,RESET);
  and AND2_2939(WX8456,WX8184,RESET);
  and AND2_2940(WX8458,WX8198,RESET);
  and AND2_2941(WX8460,WX8212,RESET);
  and AND2_2942(WX8462,WX8226,RESET);
  and AND2_2943(WX8464,WX8240,RESET);
  and AND2_2944(WX8466,WX8403,RESET);
  and AND2_2945(WX8468,WX8405,RESET);
  and AND2_2946(WX8470,WX8407,RESET);
  and AND2_2947(WX8472,WX8409,RESET);
  and AND2_2948(WX8474,WX8411,RESET);
  and AND2_2949(WX8476,WX8413,RESET);
  and AND2_2950(WX8478,WX8415,RESET);
  and AND2_2951(WX8480,WX8417,RESET);
  and AND2_2952(WX8482,WX8419,RESET);
  and AND2_2953(WX8484,WX8421,RESET);
  and AND2_2954(WX8486,WX8423,RESET);
  and AND2_2955(WX8488,WX8425,RESET);
  and AND2_2956(WX8490,WX8427,RESET);
  and AND2_2957(WX8492,WX8429,RESET);
  and AND2_2958(WX8494,WX8431,RESET);
  and AND2_2959(WX8496,WX8433,RESET);
  and AND2_2960(WX8498,WX8435,RESET);
  and AND2_2961(WX8500,WX8437,RESET);
  and AND2_2962(WX8502,WX8439,RESET);
  and AND2_2963(WX8504,WX8441,RESET);
  and AND2_2964(WX8506,WX8443,RESET);
  and AND2_2965(WX8508,WX8445,RESET);
  and AND2_2966(WX8510,WX8447,RESET);
  and AND2_2967(WX8512,WX8449,RESET);
  and AND2_2968(WX8514,WX8451,RESET);
  and AND2_2969(WX8516,WX8453,RESET);
  and AND2_2970(WX8518,WX8455,RESET);
  and AND2_2971(WX8520,WX8457,RESET);
  and AND2_2972(WX8522,WX8459,RESET);
  and AND2_2973(WX8524,WX8461,RESET);
  and AND2_2974(WX8526,WX8463,RESET);
  and AND2_2975(WX8528,WX8465,RESET);
  and AND2_2976(WX8530,WX8467,RESET);
  and AND2_2977(WX8532,WX8469,RESET);
  and AND2_2978(WX8534,WX8471,RESET);
  and AND2_2979(WX8536,WX8473,RESET);
  and AND2_2980(WX8538,WX8475,RESET);
  and AND2_2981(WX8540,WX8477,RESET);
  and AND2_2982(WX8542,WX8479,RESET);
  and AND2_2983(WX8544,WX8481,RESET);
  and AND2_2984(WX8546,WX8483,RESET);
  and AND2_2985(WX8548,WX8485,RESET);
  and AND2_2986(WX8550,WX8487,RESET);
  and AND2_2987(WX8552,WX8489,RESET);
  and AND2_2988(WX8554,WX8491,RESET);
  and AND2_2989(WX8556,WX8493,RESET);
  and AND2_2990(WX8558,WX8495,RESET);
  and AND2_2991(WX8560,WX8497,RESET);
  and AND2_2992(WX8562,WX8499,RESET);
  and AND2_2993(WX8564,WX8501,RESET);
  and AND2_2994(WX8566,WX8503,RESET);
  and AND2_2995(WX8568,WX8505,RESET);
  and AND2_2996(WX8570,WX8507,RESET);
  and AND2_2997(WX8572,WX8509,RESET);
  and AND2_2998(WX8574,WX8511,RESET);
  and AND2_2999(WX8576,WX8513,RESET);
  and AND2_3000(WX8578,WX8515,RESET);
  and AND2_3001(WX8580,WX8517,RESET);
  and AND2_3002(WX8582,WX8519,RESET);
  and AND2_3003(WX8584,WX8521,RESET);
  and AND2_3004(WX8586,WX8523,RESET);
  and AND2_3005(WX8588,WX8525,RESET);
  and AND2_3006(WX8590,WX8527,RESET);
  and AND2_3007(WX8592,WX8529,RESET);
  and AND2_3008(WX8594,WX8531,RESET);
  and AND2_3009(WX8596,WX8533,RESET);
  and AND2_3010(WX8598,WX8535,RESET);
  and AND2_3011(WX8600,WX8537,RESET);
  and AND2_3012(WX8602,WX8539,RESET);
  and AND2_3013(WX8604,WX8541,RESET);
  and AND2_3014(WX8606,WX8543,RESET);
  and AND2_3015(WX8608,WX8545,RESET);
  and AND2_3016(WX8610,WX8547,RESET);
  and AND2_3017(WX8612,WX8549,RESET);
  and AND2_3018(WX8614,WX8551,RESET);
  and AND2_3019(WX8616,WX8553,RESET);
  and AND2_3020(WX8618,WX8555,RESET);
  and AND2_3021(WX8620,WX8557,RESET);
  and AND2_3022(WX8622,WX8559,RESET);
  and AND2_3023(WX8624,WX8561,RESET);
  and AND2_3024(WX8626,WX8563,RESET);
  and AND2_3025(WX8628,WX8565,RESET);
  and AND2_3026(WX8630,WX8567,RESET);
  and AND2_3027(WX8632,WX8569,RESET);
  and AND2_3028(WX8634,WX8571,RESET);
  and AND2_3029(WX8636,WX8573,RESET);
  and AND2_3030(WX8638,WX8575,RESET);
  and AND2_3031(WX8640,WX8577,RESET);
  and AND2_3032(WX8642,WX8579,RESET);
  and AND2_3033(WX8644,WX8581,RESET);
  and AND2_3034(WX8646,WX8583,RESET);
  and AND2_3035(WX8648,WX8585,RESET);
  and AND2_3036(WX8650,WX8587,RESET);
  and AND2_3037(WX8652,WX8589,RESET);
  and AND2_3038(WX8654,WX8591,RESET);
  and AND2_3039(WX8656,WX8593,RESET);
  and AND2_3040(WX8765,WX8764,WX8763);
  and AND2_3041(WX8766,WX8338,WX8767);
  and AND2_3042(WX8772,WX8771,WX8763);
  and AND2_3043(WX8773,WX8339,WX8774);
  and AND2_3044(WX8779,WX8778,WX8763);
  and AND2_3045(WX8780,WX8340,WX8781);
  and AND2_3046(WX8786,WX8785,WX8763);
  and AND2_3047(WX8787,WX8341,WX8788);
  and AND2_3048(WX8793,WX8792,WX8763);
  and AND2_3049(WX8794,WX8342,WX8795);
  and AND2_3050(WX8800,WX8799,WX8763);
  and AND2_3051(WX8801,WX8343,WX8802);
  and AND2_3052(WX8807,WX8806,WX8763);
  and AND2_3053(WX8808,WX8344,WX8809);
  and AND2_3054(WX8814,WX8813,WX8763);
  and AND2_3055(WX8815,WX8345,WX8816);
  and AND2_3056(WX8821,WX8820,WX8763);
  and AND2_3057(WX8822,WX8346,WX8823);
  and AND2_3058(WX8828,WX8827,WX8763);
  and AND2_3059(WX8829,WX8347,WX8830);
  and AND2_3060(WX8835,WX8834,WX8763);
  and AND2_3061(WX8836,WX8348,WX8837);
  and AND2_3062(WX8842,WX8841,WX8763);
  and AND2_3063(WX8843,WX8349,WX8844);
  and AND2_3064(WX8849,WX8848,WX8763);
  and AND2_3065(WX8850,WX8350,WX8851);
  and AND2_3066(WX8856,WX8855,WX8763);
  and AND2_3067(WX8857,WX8351,WX8858);
  and AND2_3068(WX8863,WX8862,WX8763);
  and AND2_3069(WX8864,WX8352,WX8865);
  and AND2_3070(WX8870,WX8869,WX8763);
  and AND2_3071(WX8871,WX8353,WX8872);
  and AND2_3072(WX8877,WX8876,WX8763);
  and AND2_3073(WX8878,WX8354,WX8879);
  and AND2_3074(WX8884,WX8883,WX8763);
  and AND2_3075(WX8885,WX8355,WX8886);
  and AND2_3076(WX8891,WX8890,WX8763);
  and AND2_3077(WX8892,WX8356,WX8893);
  and AND2_3078(WX8898,WX8897,WX8763);
  and AND2_3079(WX8899,WX8357,WX8900);
  and AND2_3080(WX8905,WX8904,WX8763);
  and AND2_3081(WX8906,WX8358,WX8907);
  and AND2_3082(WX8912,WX8911,WX8763);
  and AND2_3083(WX8913,WX8359,WX8914);
  and AND2_3084(WX8919,WX8918,WX8763);
  and AND2_3085(WX8920,WX8360,WX8921);
  and AND2_3086(WX8926,WX8925,WX8763);
  and AND2_3087(WX8927,WX8361,WX8928);
  and AND2_3088(WX8933,WX8932,WX8763);
  and AND2_3089(WX8934,WX8362,WX8935);
  and AND2_3090(WX8940,WX8939,WX8763);
  and AND2_3091(WX8941,WX8363,WX8942);
  and AND2_3092(WX8947,WX8946,WX8763);
  and AND2_3093(WX8948,WX8364,WX8949);
  and AND2_3094(WX8954,WX8953,WX8763);
  and AND2_3095(WX8955,WX8365,WX8956);
  and AND2_3096(WX8961,WX8960,WX8763);
  and AND2_3097(WX8962,WX8366,WX8963);
  and AND2_3098(WX8968,WX8967,WX8763);
  and AND2_3099(WX8969,WX8367,WX8970);
  and AND2_3100(WX8975,WX8974,WX8763);
  and AND2_3101(WX8976,WX8368,WX8977);
  and AND2_3102(WX8982,WX8981,WX8763);
  and AND2_3103(WX8983,WX8369,WX8984);
  and AND2_3104(WX9022,WX8992,WX9021);
  and AND2_3105(WX9024,WX9020,WX9021);
  and AND2_3106(WX9026,WX9019,WX9021);
  and AND2_3107(WX9028,WX9018,WX9021);
  and AND2_3108(WX9030,WX8991,WX9021);
  and AND2_3109(WX9032,WX9017,WX9021);
  and AND2_3110(WX9034,WX9016,WX9021);
  and AND2_3111(WX9036,WX9015,WX9021);
  and AND2_3112(WX9038,WX9014,WX9021);
  and AND2_3113(WX9040,WX9013,WX9021);
  and AND2_3114(WX9042,WX9012,WX9021);
  and AND2_3115(WX9044,WX8990,WX9021);
  and AND2_3116(WX9046,WX9011,WX9021);
  and AND2_3117(WX9048,WX9010,WX9021);
  and AND2_3118(WX9050,WX9009,WX9021);
  and AND2_3119(WX9052,WX9008,WX9021);
  and AND2_3120(WX9054,WX8989,WX9021);
  and AND2_3121(WX9056,WX9007,WX9021);
  and AND2_3122(WX9058,WX9006,WX9021);
  and AND2_3123(WX9060,WX9005,WX9021);
  and AND2_3124(WX9062,WX9004,WX9021);
  and AND2_3125(WX9064,WX9003,WX9021);
  and AND2_3126(WX9066,WX9002,WX9021);
  and AND2_3127(WX9068,WX9001,WX9021);
  and AND2_3128(WX9070,WX9000,WX9021);
  and AND2_3129(WX9072,WX8999,WX9021);
  and AND2_3130(WX9074,WX8998,WX9021);
  and AND2_3131(WX9076,WX8997,WX9021);
  and AND2_3132(WX9078,WX8996,WX9021);
  and AND2_3133(WX9080,WX8995,WX9021);
  and AND2_3134(WX9082,WX8994,WX9021);
  and AND2_3135(WX9084,WX8993,WX9021);
  and AND2_3136(WX9086,WX9097,WX10054);
  and AND2_3137(WX9087,WX9093,WX9088);
  and AND2_3138(WX9090,CRC_OUT_2_31,WX10055);
  and AND2_3139(WX9091,WX11356,WX9092);
  and AND2_3140(WX9094,WX9536,WX10055);
  and AND2_3141(WX9095,WX10063,WX9096);
  and AND2_3142(WX9100,WX9111,WX10054);
  and AND2_3143(WX9101,WX9107,WX9102);
  and AND2_3144(WX9104,CRC_OUT_2_30,WX10055);
  and AND2_3145(WX9105,WX11363,WX9106);
  and AND2_3146(WX9108,WX9538,WX10055);
  and AND2_3147(WX9109,WX10070,WX9110);
  and AND2_3148(WX9114,WX9125,WX10054);
  and AND2_3149(WX9115,WX9121,WX9116);
  and AND2_3150(WX9118,CRC_OUT_2_29,WX10055);
  and AND2_3151(WX9119,WX11370,WX9120);
  and AND2_3152(WX9122,WX9540,WX10055);
  and AND2_3153(WX9123,WX10077,WX9124);
  and AND2_3154(WX9128,WX9139,WX10054);
  and AND2_3155(WX9129,WX9135,WX9130);
  and AND2_3156(WX9132,CRC_OUT_2_28,WX10055);
  and AND2_3157(WX9133,WX11377,WX9134);
  and AND2_3158(WX9136,WX9542,WX10055);
  and AND2_3159(WX9137,WX10084,WX9138);
  and AND2_3160(WX9142,WX9153,WX10054);
  and AND2_3161(WX9143,WX9149,WX9144);
  and AND2_3162(WX9146,CRC_OUT_2_27,WX10055);
  and AND2_3163(WX9147,WX11384,WX9148);
  and AND2_3164(WX9150,WX9544,WX10055);
  and AND2_3165(WX9151,WX10091,WX9152);
  and AND2_3166(WX9156,WX9167,WX10054);
  and AND2_3167(WX9157,WX9163,WX9158);
  and AND2_3168(WX9160,CRC_OUT_2_26,WX10055);
  and AND2_3169(WX9161,WX11391,WX9162);
  and AND2_3170(WX9164,WX9546,WX10055);
  and AND2_3171(WX9165,WX10098,WX9166);
  and AND2_3172(WX9170,WX9181,WX10054);
  and AND2_3173(WX9171,WX9177,WX9172);
  and AND2_3174(WX9174,CRC_OUT_2_25,WX10055);
  and AND2_3175(WX9175,WX11398,WX9176);
  and AND2_3176(WX9178,WX9548,WX10055);
  and AND2_3177(WX9179,WX10105,WX9180);
  and AND2_3178(WX9184,WX9195,WX10054);
  and AND2_3179(WX9185,WX9191,WX9186);
  and AND2_3180(WX9188,CRC_OUT_2_24,WX10055);
  and AND2_3181(WX9189,WX11405,WX9190);
  and AND2_3182(WX9192,WX9550,WX10055);
  and AND2_3183(WX9193,WX10112,WX9194);
  and AND2_3184(WX9198,WX9209,WX10054);
  and AND2_3185(WX9199,WX9205,WX9200);
  and AND2_3186(WX9202,CRC_OUT_2_23,WX10055);
  and AND2_3187(WX9203,WX11412,WX9204);
  and AND2_3188(WX9206,WX9552,WX10055);
  and AND2_3189(WX9207,WX10119,WX9208);
  and AND2_3190(WX9212,WX9223,WX10054);
  and AND2_3191(WX9213,WX9219,WX9214);
  and AND2_3192(WX9216,CRC_OUT_2_22,WX10055);
  and AND2_3193(WX9217,WX11419,WX9218);
  and AND2_3194(WX9220,WX9554,WX10055);
  and AND2_3195(WX9221,WX10126,WX9222);
  and AND2_3196(WX9226,WX9237,WX10054);
  and AND2_3197(WX9227,WX9233,WX9228);
  and AND2_3198(WX9230,CRC_OUT_2_21,WX10055);
  and AND2_3199(WX9231,WX11426,WX9232);
  and AND2_3200(WX9234,WX9556,WX10055);
  and AND2_3201(WX9235,WX10133,WX9236);
  and AND2_3202(WX9240,WX9251,WX10054);
  and AND2_3203(WX9241,WX9247,WX9242);
  and AND2_3204(WX9244,CRC_OUT_2_20,WX10055);
  and AND2_3205(WX9245,WX11433,WX9246);
  and AND2_3206(WX9248,WX9558,WX10055);
  and AND2_3207(WX9249,WX10140,WX9250);
  and AND2_3208(WX9254,WX9265,WX10054);
  and AND2_3209(WX9255,WX9261,WX9256);
  and AND2_3210(WX9258,CRC_OUT_2_19,WX10055);
  and AND2_3211(WX9259,WX11440,WX9260);
  and AND2_3212(WX9262,WX9560,WX10055);
  and AND2_3213(WX9263,WX10147,WX9264);
  and AND2_3214(WX9268,WX9279,WX10054);
  and AND2_3215(WX9269,WX9275,WX9270);
  and AND2_3216(WX9272,CRC_OUT_2_18,WX10055);
  and AND2_3217(WX9273,WX11447,WX9274);
  and AND2_3218(WX9276,WX9562,WX10055);
  and AND2_3219(WX9277,WX10154,WX9278);
  and AND2_3220(WX9282,WX9293,WX10054);
  and AND2_3221(WX9283,WX9289,WX9284);
  and AND2_3222(WX9286,CRC_OUT_2_17,WX10055);
  and AND2_3223(WX9287,WX11454,WX9288);
  and AND2_3224(WX9290,WX9564,WX10055);
  and AND2_3225(WX9291,WX10161,WX9292);
  and AND2_3226(WX9296,WX9307,WX10054);
  and AND2_3227(WX9297,WX9303,WX9298);
  and AND2_3228(WX9300,CRC_OUT_2_16,WX10055);
  and AND2_3229(WX9301,WX11461,WX9302);
  and AND2_3230(WX9304,WX9566,WX10055);
  and AND2_3231(WX9305,WX10168,WX9306);
  and AND2_3232(WX9310,WX9321,WX10054);
  and AND2_3233(WX9311,WX9317,WX9312);
  and AND2_3234(WX9314,CRC_OUT_2_15,WX10055);
  and AND2_3235(WX9315,WX11468,WX9316);
  and AND2_3236(WX9318,WX9568,WX10055);
  and AND2_3237(WX9319,WX10175,WX9320);
  and AND2_3238(WX9324,WX9335,WX10054);
  and AND2_3239(WX9325,WX9331,WX9326);
  and AND2_3240(WX9328,CRC_OUT_2_14,WX10055);
  and AND2_3241(WX9329,WX11475,WX9330);
  and AND2_3242(WX9332,WX9570,WX10055);
  and AND2_3243(WX9333,WX10182,WX9334);
  and AND2_3244(WX9338,WX9349,WX10054);
  and AND2_3245(WX9339,WX9345,WX9340);
  and AND2_3246(WX9342,CRC_OUT_2_13,WX10055);
  and AND2_3247(WX9343,WX11482,WX9344);
  and AND2_3248(WX9346,WX9572,WX10055);
  and AND2_3249(WX9347,WX10189,WX9348);
  and AND2_3250(WX9352,WX9363,WX10054);
  and AND2_3251(WX9353,WX9359,WX9354);
  and AND2_3252(WX9356,CRC_OUT_2_12,WX10055);
  and AND2_3253(WX9357,WX11489,WX9358);
  and AND2_3254(WX9360,WX9574,WX10055);
  and AND2_3255(WX9361,WX10196,WX9362);
  and AND2_3256(WX9366,WX9377,WX10054);
  and AND2_3257(WX9367,WX9373,WX9368);
  and AND2_3258(WX9370,CRC_OUT_2_11,WX10055);
  and AND2_3259(WX9371,WX11496,WX9372);
  and AND2_3260(WX9374,WX9576,WX10055);
  and AND2_3261(WX9375,WX10203,WX9376);
  and AND2_3262(WX9380,WX9391,WX10054);
  and AND2_3263(WX9381,WX9387,WX9382);
  and AND2_3264(WX9384,CRC_OUT_2_10,WX10055);
  and AND2_3265(WX9385,WX11503,WX9386);
  and AND2_3266(WX9388,WX9578,WX10055);
  and AND2_3267(WX9389,WX10210,WX9390);
  and AND2_3268(WX9394,WX9405,WX10054);
  and AND2_3269(WX9395,WX9401,WX9396);
  and AND2_3270(WX9398,CRC_OUT_2_9,WX10055);
  and AND2_3271(WX9399,WX11510,WX9400);
  and AND2_3272(WX9402,WX9580,WX10055);
  and AND2_3273(WX9403,WX10217,WX9404);
  and AND2_3274(WX9408,WX9419,WX10054);
  and AND2_3275(WX9409,WX9415,WX9410);
  and AND2_3276(WX9412,CRC_OUT_2_8,WX10055);
  and AND2_3277(WX9413,WX11517,WX9414);
  and AND2_3278(WX9416,WX9582,WX10055);
  and AND2_3279(WX9417,WX10224,WX9418);
  and AND2_3280(WX9422,WX9433,WX10054);
  and AND2_3281(WX9423,WX9429,WX9424);
  and AND2_3282(WX9426,CRC_OUT_2_7,WX10055);
  and AND2_3283(WX9427,WX11524,WX9428);
  and AND2_3284(WX9430,WX9584,WX10055);
  and AND2_3285(WX9431,WX10231,WX9432);
  and AND2_3286(WX9436,WX9447,WX10054);
  and AND2_3287(WX9437,WX9443,WX9438);
  and AND2_3288(WX9440,CRC_OUT_2_6,WX10055);
  and AND2_3289(WX9441,WX11531,WX9442);
  and AND2_3290(WX9444,WX9586,WX10055);
  and AND2_3291(WX9445,WX10238,WX9446);
  and AND2_3292(WX9450,WX9461,WX10054);
  and AND2_3293(WX9451,WX9457,WX9452);
  and AND2_3294(WX9454,CRC_OUT_2_5,WX10055);
  and AND2_3295(WX9455,WX11538,WX9456);
  and AND2_3296(WX9458,WX9588,WX10055);
  and AND2_3297(WX9459,WX10245,WX9460);
  and AND2_3298(WX9464,WX9475,WX10054);
  and AND2_3299(WX9465,WX9471,WX9466);
  and AND2_3300(WX9468,CRC_OUT_2_4,WX10055);
  and AND2_3301(WX9469,WX11545,WX9470);
  and AND2_3302(WX9472,WX9590,WX10055);
  and AND2_3303(WX9473,WX10252,WX9474);
  and AND2_3304(WX9478,WX9489,WX10054);
  and AND2_3305(WX9479,WX9485,WX9480);
  and AND2_3306(WX9482,CRC_OUT_2_3,WX10055);
  and AND2_3307(WX9483,WX11552,WX9484);
  and AND2_3308(WX9486,WX9592,WX10055);
  and AND2_3309(WX9487,WX10259,WX9488);
  and AND2_3310(WX9492,WX9503,WX10054);
  and AND2_3311(WX9493,WX9499,WX9494);
  and AND2_3312(WX9496,CRC_OUT_2_2,WX10055);
  and AND2_3313(WX9497,WX11559,WX9498);
  and AND2_3314(WX9500,WX9594,WX10055);
  and AND2_3315(WX9501,WX10266,WX9502);
  and AND2_3316(WX9506,WX9517,WX10054);
  and AND2_3317(WX9507,WX9513,WX9508);
  and AND2_3318(WX9510,CRC_OUT_2_1,WX10055);
  and AND2_3319(WX9511,WX11566,WX9512);
  and AND2_3320(WX9514,WX9596,WX10055);
  and AND2_3321(WX9515,WX10273,WX9516);
  and AND2_3322(WX9520,WX9531,WX10054);
  and AND2_3323(WX9521,WX9527,WX9522);
  and AND2_3324(WX9524,CRC_OUT_2_0,WX10055);
  and AND2_3325(WX9525,WX11573,WX9526);
  and AND2_3326(WX9528,WX9598,WX10055);
  and AND2_3327(WX9529,WX10280,WX9530);
  and AND2_3328(WX9535,WX9538,RESET);
  and AND2_3329(WX9537,WX9540,RESET);
  and AND2_3330(WX9539,WX9542,RESET);
  and AND2_3331(WX9541,WX9544,RESET);
  and AND2_3332(WX9543,WX9546,RESET);
  and AND2_3333(WX9545,WX9548,RESET);
  and AND2_3334(WX9547,WX9550,RESET);
  and AND2_3335(WX9549,WX9552,RESET);
  and AND2_3336(WX9551,WX9554,RESET);
  and AND2_3337(WX9553,WX9556,RESET);
  and AND2_3338(WX9555,WX9558,RESET);
  and AND2_3339(WX9557,WX9560,RESET);
  and AND2_3340(WX9559,WX9562,RESET);
  and AND2_3341(WX9561,WX9564,RESET);
  and AND2_3342(WX9563,WX9566,RESET);
  and AND2_3343(WX9565,WX9568,RESET);
  and AND2_3344(WX9567,WX9570,RESET);
  and AND2_3345(WX9569,WX9572,RESET);
  and AND2_3346(WX9571,WX9574,RESET);
  and AND2_3347(WX9573,WX9576,RESET);
  and AND2_3348(WX9575,WX9578,RESET);
  and AND2_3349(WX9577,WX9580,RESET);
  and AND2_3350(WX9579,WX9582,RESET);
  and AND2_3351(WX9581,WX9584,RESET);
  and AND2_3352(WX9583,WX9586,RESET);
  and AND2_3353(WX9585,WX9588,RESET);
  and AND2_3354(WX9587,WX9590,RESET);
  and AND2_3355(WX9589,WX9592,RESET);
  and AND2_3356(WX9591,WX9594,RESET);
  and AND2_3357(WX9593,WX9596,RESET);
  and AND2_3358(WX9595,WX9598,RESET);
  and AND2_3359(WX9597,WX9534,RESET);
  and AND2_3360(WX9695,WX9099,RESET);
  and AND2_3361(WX9697,WX9113,RESET);
  and AND2_3362(WX9699,WX9127,RESET);
  and AND2_3363(WX9701,WX9141,RESET);
  and AND2_3364(WX9703,WX9155,RESET);
  and AND2_3365(WX9705,WX9169,RESET);
  and AND2_3366(WX9707,WX9183,RESET);
  and AND2_3367(WX9709,WX9197,RESET);
  and AND2_3368(WX9711,WX9211,RESET);
  and AND2_3369(WX9713,WX9225,RESET);
  and AND2_3370(WX9715,WX9239,RESET);
  and AND2_3371(WX9717,WX9253,RESET);
  and AND2_3372(WX9719,WX9267,RESET);
  and AND2_3373(WX9721,WX9281,RESET);
  and AND2_3374(WX9723,WX9295,RESET);
  and AND2_3375(WX9725,WX9309,RESET);
  and AND2_3376(WX9727,WX9323,RESET);
  and AND2_3377(WX9729,WX9337,RESET);
  and AND2_3378(WX9731,WX9351,RESET);
  and AND2_3379(WX9733,WX9365,RESET);
  and AND2_3380(WX9735,WX9379,RESET);
  and AND2_3381(WX9737,WX9393,RESET);
  and AND2_3382(WX9739,WX9407,RESET);
  and AND2_3383(WX9741,WX9421,RESET);
  and AND2_3384(WX9743,WX9435,RESET);
  and AND2_3385(WX9745,WX9449,RESET);
  and AND2_3386(WX9747,WX9463,RESET);
  and AND2_3387(WX9749,WX9477,RESET);
  and AND2_3388(WX9751,WX9491,RESET);
  and AND2_3389(WX9753,WX9505,RESET);
  and AND2_3390(WX9755,WX9519,RESET);
  and AND2_3391(WX9757,WX9533,RESET);
  and AND2_3392(WX9759,WX9696,RESET);
  and AND2_3393(WX9761,WX9698,RESET);
  and AND2_3394(WX9763,WX9700,RESET);
  and AND2_3395(WX9765,WX9702,RESET);
  and AND2_3396(WX9767,WX9704,RESET);
  and AND2_3397(WX9769,WX9706,RESET);
  and AND2_3398(WX9771,WX9708,RESET);
  and AND2_3399(WX9773,WX9710,RESET);
  and AND2_3400(WX9775,WX9712,RESET);
  and AND2_3401(WX9777,WX9714,RESET);
  and AND2_3402(WX9779,WX9716,RESET);
  and AND2_3403(WX9781,WX9718,RESET);
  and AND2_3404(WX9783,WX9720,RESET);
  and AND2_3405(WX9785,WX9722,RESET);
  and AND2_3406(WX9787,WX9724,RESET);
  and AND2_3407(WX9789,WX9726,RESET);
  and AND2_3408(WX9791,WX9728,RESET);
  and AND2_3409(WX9793,WX9730,RESET);
  and AND2_3410(WX9795,WX9732,RESET);
  and AND2_3411(WX9797,WX9734,RESET);
  and AND2_3412(WX9799,WX9736,RESET);
  and AND2_3413(WX9801,WX9738,RESET);
  and AND2_3414(WX9803,WX9740,RESET);
  and AND2_3415(WX9805,WX9742,RESET);
  and AND2_3416(WX9807,WX9744,RESET);
  and AND2_3417(WX9809,WX9746,RESET);
  and AND2_3418(WX9811,WX9748,RESET);
  and AND2_3419(WX9813,WX9750,RESET);
  and AND2_3420(WX9815,WX9752,RESET);
  and AND2_3421(WX9817,WX9754,RESET);
  and AND2_3422(WX9819,WX9756,RESET);
  and AND2_3423(WX9821,WX9758,RESET);
  and AND2_3424(WX9823,WX9760,RESET);
  and AND2_3425(WX9825,WX9762,RESET);
  and AND2_3426(WX9827,WX9764,RESET);
  and AND2_3427(WX9829,WX9766,RESET);
  and AND2_3428(WX9831,WX9768,RESET);
  and AND2_3429(WX9833,WX9770,RESET);
  and AND2_3430(WX9835,WX9772,RESET);
  and AND2_3431(WX9837,WX9774,RESET);
  and AND2_3432(WX9839,WX9776,RESET);
  and AND2_3433(WX9841,WX9778,RESET);
  and AND2_3434(WX9843,WX9780,RESET);
  and AND2_3435(WX9845,WX9782,RESET);
  and AND2_3436(WX9847,WX9784,RESET);
  and AND2_3437(WX9849,WX9786,RESET);
  and AND2_3438(WX9851,WX9788,RESET);
  and AND2_3439(WX9853,WX9790,RESET);
  and AND2_3440(WX9855,WX9792,RESET);
  and AND2_3441(WX9857,WX9794,RESET);
  and AND2_3442(WX9859,WX9796,RESET);
  and AND2_3443(WX9861,WX9798,RESET);
  and AND2_3444(WX9863,WX9800,RESET);
  and AND2_3445(WX9865,WX9802,RESET);
  and AND2_3446(WX9867,WX9804,RESET);
  and AND2_3447(WX9869,WX9806,RESET);
  and AND2_3448(WX9871,WX9808,RESET);
  and AND2_3449(WX9873,WX9810,RESET);
  and AND2_3450(WX9875,WX9812,RESET);
  and AND2_3451(WX9877,WX9814,RESET);
  and AND2_3452(WX9879,WX9816,RESET);
  and AND2_3453(WX9881,WX9818,RESET);
  and AND2_3454(WX9883,WX9820,RESET);
  and AND2_3455(WX9885,WX9822,RESET);
  and AND2_3456(WX9887,WX9824,RESET);
  and AND2_3457(WX9889,WX9826,RESET);
  and AND2_3458(WX9891,WX9828,RESET);
  and AND2_3459(WX9893,WX9830,RESET);
  and AND2_3460(WX9895,WX9832,RESET);
  and AND2_3461(WX9897,WX9834,RESET);
  and AND2_3462(WX9899,WX9836,RESET);
  and AND2_3463(WX9901,WX9838,RESET);
  and AND2_3464(WX9903,WX9840,RESET);
  and AND2_3465(WX9905,WX9842,RESET);
  and AND2_3466(WX9907,WX9844,RESET);
  and AND2_3467(WX9909,WX9846,RESET);
  and AND2_3468(WX9911,WX9848,RESET);
  and AND2_3469(WX9913,WX9850,RESET);
  and AND2_3470(WX9915,WX9852,RESET);
  and AND2_3471(WX9917,WX9854,RESET);
  and AND2_3472(WX9919,WX9856,RESET);
  and AND2_3473(WX9921,WX9858,RESET);
  and AND2_3474(WX9923,WX9860,RESET);
  and AND2_3475(WX9925,WX9862,RESET);
  and AND2_3476(WX9927,WX9864,RESET);
  and AND2_3477(WX9929,WX9866,RESET);
  and AND2_3478(WX9931,WX9868,RESET);
  and AND2_3479(WX9933,WX9870,RESET);
  and AND2_3480(WX9935,WX9872,RESET);
  and AND2_3481(WX9937,WX9874,RESET);
  and AND2_3482(WX9939,WX9876,RESET);
  and AND2_3483(WX9941,WX9878,RESET);
  and AND2_3484(WX9943,WX9880,RESET);
  and AND2_3485(WX9945,WX9882,RESET);
  and AND2_3486(WX9947,WX9884,RESET);
  and AND2_3487(WX9949,WX9886,RESET);
  and AND2_3488(WX10058,WX10057,WX10056);
  and AND2_3489(WX10059,WX9631,WX10060);
  and AND2_3490(WX10065,WX10064,WX10056);
  and AND2_3491(WX10066,WX9632,WX10067);
  and AND2_3492(WX10072,WX10071,WX10056);
  and AND2_3493(WX10073,WX9633,WX10074);
  and AND2_3494(WX10079,WX10078,WX10056);
  and AND2_3495(WX10080,WX9634,WX10081);
  and AND2_3496(WX10086,WX10085,WX10056);
  and AND2_3497(WX10087,WX9635,WX10088);
  and AND2_3498(WX10093,WX10092,WX10056);
  and AND2_3499(WX10094,WX9636,WX10095);
  and AND2_3500(WX10100,WX10099,WX10056);
  and AND2_3501(WX10101,WX9637,WX10102);
  and AND2_3502(WX10107,WX10106,WX10056);
  and AND2_3503(WX10108,WX9638,WX10109);
  and AND2_3504(WX10114,WX10113,WX10056);
  and AND2_3505(WX10115,WX9639,WX10116);
  and AND2_3506(WX10121,WX10120,WX10056);
  and AND2_3507(WX10122,WX9640,WX10123);
  and AND2_3508(WX10128,WX10127,WX10056);
  and AND2_3509(WX10129,WX9641,WX10130);
  and AND2_3510(WX10135,WX10134,WX10056);
  and AND2_3511(WX10136,WX9642,WX10137);
  and AND2_3512(WX10142,WX10141,WX10056);
  and AND2_3513(WX10143,WX9643,WX10144);
  and AND2_3514(WX10149,WX10148,WX10056);
  and AND2_3515(WX10150,WX9644,WX10151);
  and AND2_3516(WX10156,WX10155,WX10056);
  and AND2_3517(WX10157,WX9645,WX10158);
  and AND2_3518(WX10163,WX10162,WX10056);
  and AND2_3519(WX10164,WX9646,WX10165);
  and AND2_3520(WX10170,WX10169,WX10056);
  and AND2_3521(WX10171,WX9647,WX10172);
  and AND2_3522(WX10177,WX10176,WX10056);
  and AND2_3523(WX10178,WX9648,WX10179);
  and AND2_3524(WX10184,WX10183,WX10056);
  and AND2_3525(WX10185,WX9649,WX10186);
  and AND2_3526(WX10191,WX10190,WX10056);
  and AND2_3527(WX10192,WX9650,WX10193);
  and AND2_3528(WX10198,WX10197,WX10056);
  and AND2_3529(WX10199,WX9651,WX10200);
  and AND2_3530(WX10205,WX10204,WX10056);
  and AND2_3531(WX10206,WX9652,WX10207);
  and AND2_3532(WX10212,WX10211,WX10056);
  and AND2_3533(WX10213,WX9653,WX10214);
  and AND2_3534(WX10219,WX10218,WX10056);
  and AND2_3535(WX10220,WX9654,WX10221);
  and AND2_3536(WX10226,WX10225,WX10056);
  and AND2_3537(WX10227,WX9655,WX10228);
  and AND2_3538(WX10233,WX10232,WX10056);
  and AND2_3539(WX10234,WX9656,WX10235);
  and AND2_3540(WX10240,WX10239,WX10056);
  and AND2_3541(WX10241,WX9657,WX10242);
  and AND2_3542(WX10247,WX10246,WX10056);
  and AND2_3543(WX10248,WX9658,WX10249);
  and AND2_3544(WX10254,WX10253,WX10056);
  and AND2_3545(WX10255,WX9659,WX10256);
  and AND2_3546(WX10261,WX10260,WX10056);
  and AND2_3547(WX10262,WX9660,WX10263);
  and AND2_3548(WX10268,WX10267,WX10056);
  and AND2_3549(WX10269,WX9661,WX10270);
  and AND2_3550(WX10275,WX10274,WX10056);
  and AND2_3551(WX10276,WX9662,WX10277);
  and AND2_3552(WX10315,WX10285,WX10314);
  and AND2_3553(WX10317,WX10313,WX10314);
  and AND2_3554(WX10319,WX10312,WX10314);
  and AND2_3555(WX10321,WX10311,WX10314);
  and AND2_3556(WX10323,WX10284,WX10314);
  and AND2_3557(WX10325,WX10310,WX10314);
  and AND2_3558(WX10327,WX10309,WX10314);
  and AND2_3559(WX10329,WX10308,WX10314);
  and AND2_3560(WX10331,WX10307,WX10314);
  and AND2_3561(WX10333,WX10306,WX10314);
  and AND2_3562(WX10335,WX10305,WX10314);
  and AND2_3563(WX10337,WX10283,WX10314);
  and AND2_3564(WX10339,WX10304,WX10314);
  and AND2_3565(WX10341,WX10303,WX10314);
  and AND2_3566(WX10343,WX10302,WX10314);
  and AND2_3567(WX10345,WX10301,WX10314);
  and AND2_3568(WX10347,WX10282,WX10314);
  and AND2_3569(WX10349,WX10300,WX10314);
  and AND2_3570(WX10351,WX10299,WX10314);
  and AND2_3571(WX10353,WX10298,WX10314);
  and AND2_3572(WX10355,WX10297,WX10314);
  and AND2_3573(WX10357,WX10296,WX10314);
  and AND2_3574(WX10359,WX10295,WX10314);
  and AND2_3575(WX10361,WX10294,WX10314);
  and AND2_3576(WX10363,WX10293,WX10314);
  and AND2_3577(WX10365,WX10292,WX10314);
  and AND2_3578(WX10367,WX10291,WX10314);
  and AND2_3579(WX10369,WX10290,WX10314);
  and AND2_3580(WX10371,WX10289,WX10314);
  and AND2_3581(WX10373,WX10288,WX10314);
  and AND2_3582(WX10375,WX10287,WX10314);
  and AND2_3583(WX10377,WX10286,WX10314);
  and AND2_3584(WX10379,WX10390,WX11347);
  and AND2_3585(WX10380,WX10386,WX10381);
  and AND2_3586(WX10383,CRC_OUT_1_31,WX11348);
  and AND2_3587(WX10384,DATA_0_31,WX10385);
  and AND2_3588(WX10387,WX10829,WX11348);
  and AND2_3589(WX10388,WX11356,WX10389);
  and AND2_3590(WX10393,WX10404,WX11347);
  and AND2_3591(WX10394,WX10400,WX10395);
  and AND2_3592(WX10397,CRC_OUT_1_30,WX11348);
  and AND2_3593(WX10398,DATA_0_30,WX10399);
  and AND2_3594(WX10401,WX10831,WX11348);
  and AND2_3595(WX10402,WX11363,WX10403);
  and AND2_3596(WX10407,WX10418,WX11347);
  and AND2_3597(WX10408,WX10414,WX10409);
  and AND2_3598(WX10411,CRC_OUT_1_29,WX11348);
  and AND2_3599(WX10412,DATA_0_29,WX10413);
  and AND2_3600(WX10415,WX10833,WX11348);
  and AND2_3601(WX10416,WX11370,WX10417);
  and AND2_3602(WX10421,WX10432,WX11347);
  and AND2_3603(WX10422,WX10428,WX10423);
  and AND2_3604(WX10425,CRC_OUT_1_28,WX11348);
  and AND2_3605(WX10426,DATA_0_28,WX10427);
  and AND2_3606(WX10429,WX10835,WX11348);
  and AND2_3607(WX10430,WX11377,WX10431);
  and AND2_3608(WX10435,WX10446,WX11347);
  and AND2_3609(WX10436,WX10442,WX10437);
  and AND2_3610(WX10439,CRC_OUT_1_27,WX11348);
  and AND2_3611(WX10440,DATA_0_27,WX10441);
  and AND2_3612(WX10443,WX10837,WX11348);
  and AND2_3613(WX10444,WX11384,WX10445);
  and AND2_3614(WX10449,WX10460,WX11347);
  and AND2_3615(WX10450,WX10456,WX10451);
  and AND2_3616(WX10453,CRC_OUT_1_26,WX11348);
  and AND2_3617(WX10454,DATA_0_26,WX10455);
  and AND2_3618(WX10457,WX10839,WX11348);
  and AND2_3619(WX10458,WX11391,WX10459);
  and AND2_3620(WX10463,WX10474,WX11347);
  and AND2_3621(WX10464,WX10470,WX10465);
  and AND2_3622(WX10467,CRC_OUT_1_25,WX11348);
  and AND2_3623(WX10468,DATA_0_25,WX10469);
  and AND2_3624(WX10471,WX10841,WX11348);
  and AND2_3625(WX10472,WX11398,WX10473);
  and AND2_3626(WX10477,WX10488,WX11347);
  and AND2_3627(WX10478,WX10484,WX10479);
  and AND2_3628(WX10481,CRC_OUT_1_24,WX11348);
  and AND2_3629(WX10482,DATA_0_24,WX10483);
  and AND2_3630(WX10485,WX10843,WX11348);
  and AND2_3631(WX10486,WX11405,WX10487);
  and AND2_3632(WX10491,WX10502,WX11347);
  and AND2_3633(WX10492,WX10498,WX10493);
  and AND2_3634(WX10495,CRC_OUT_1_23,WX11348);
  and AND2_3635(WX10496,DATA_0_23,WX10497);
  and AND2_3636(WX10499,WX10845,WX11348);
  and AND2_3637(WX10500,WX11412,WX10501);
  and AND2_3638(WX10505,WX10516,WX11347);
  and AND2_3639(WX10506,WX10512,WX10507);
  and AND2_3640(WX10509,CRC_OUT_1_22,WX11348);
  and AND2_3641(WX10510,DATA_0_22,WX10511);
  and AND2_3642(WX10513,WX10847,WX11348);
  and AND2_3643(WX10514,WX11419,WX10515);
  and AND2_3644(WX10519,WX10530,WX11347);
  and AND2_3645(WX10520,WX10526,WX10521);
  and AND2_3646(WX10523,CRC_OUT_1_21,WX11348);
  and AND2_3647(WX10524,DATA_0_21,WX10525);
  and AND2_3648(WX10527,WX10849,WX11348);
  and AND2_3649(WX10528,WX11426,WX10529);
  and AND2_3650(WX10533,WX10544,WX11347);
  and AND2_3651(WX10534,WX10540,WX10535);
  and AND2_3652(WX10537,CRC_OUT_1_20,WX11348);
  and AND2_3653(WX10538,DATA_0_20,WX10539);
  and AND2_3654(WX10541,WX10851,WX11348);
  and AND2_3655(WX10542,WX11433,WX10543);
  and AND2_3656(WX10547,WX10558,WX11347);
  and AND2_3657(WX10548,WX10554,WX10549);
  and AND2_3658(WX10551,CRC_OUT_1_19,WX11348);
  and AND2_3659(WX10552,DATA_0_19,WX10553);
  and AND2_3660(WX10555,WX10853,WX11348);
  and AND2_3661(WX10556,WX11440,WX10557);
  and AND2_3662(WX10561,WX10572,WX11347);
  and AND2_3663(WX10562,WX10568,WX10563);
  and AND2_3664(WX10565,CRC_OUT_1_18,WX11348);
  and AND2_3665(WX10566,DATA_0_18,WX10567);
  and AND2_3666(WX10569,WX10855,WX11348);
  and AND2_3667(WX10570,WX11447,WX10571);
  and AND2_3668(WX10575,WX10586,WX11347);
  and AND2_3669(WX10576,WX10582,WX10577);
  and AND2_3670(WX10579,CRC_OUT_1_17,WX11348);
  and AND2_3671(WX10580,DATA_0_17,WX10581);
  and AND2_3672(WX10583,WX10857,WX11348);
  and AND2_3673(WX10584,WX11454,WX10585);
  and AND2_3674(WX10589,WX10600,WX11347);
  and AND2_3675(WX10590,WX10596,WX10591);
  and AND2_3676(WX10593,CRC_OUT_1_16,WX11348);
  and AND2_3677(WX10594,DATA_0_16,WX10595);
  and AND2_3678(WX10597,WX10859,WX11348);
  and AND2_3679(WX10598,WX11461,WX10599);
  and AND2_3680(WX10603,WX10614,WX11347);
  and AND2_3681(WX10604,WX10610,WX10605);
  and AND2_3682(WX10607,CRC_OUT_1_15,WX11348);
  and AND2_3683(WX10608,DATA_0_15,WX10609);
  and AND2_3684(WX10611,WX10861,WX11348);
  and AND2_3685(WX10612,WX11468,WX10613);
  and AND2_3686(WX10617,WX10628,WX11347);
  and AND2_3687(WX10618,WX10624,WX10619);
  and AND2_3688(WX10621,CRC_OUT_1_14,WX11348);
  and AND2_3689(WX10622,DATA_0_14,WX10623);
  and AND2_3690(WX10625,WX10863,WX11348);
  and AND2_3691(WX10626,WX11475,WX10627);
  and AND2_3692(WX10631,WX10642,WX11347);
  and AND2_3693(WX10632,WX10638,WX10633);
  and AND2_3694(WX10635,CRC_OUT_1_13,WX11348);
  and AND2_3695(WX10636,DATA_0_13,WX10637);
  and AND2_3696(WX10639,WX10865,WX11348);
  and AND2_3697(WX10640,WX11482,WX10641);
  and AND2_3698(WX10645,WX10656,WX11347);
  and AND2_3699(WX10646,WX10652,WX10647);
  and AND2_3700(WX10649,CRC_OUT_1_12,WX11348);
  and AND2_3701(WX10650,DATA_0_12,WX10651);
  and AND2_3702(WX10653,WX10867,WX11348);
  and AND2_3703(WX10654,WX11489,WX10655);
  and AND2_3704(WX10659,WX10670,WX11347);
  and AND2_3705(WX10660,WX10666,WX10661);
  and AND2_3706(WX10663,CRC_OUT_1_11,WX11348);
  and AND2_3707(WX10664,DATA_0_11,WX10665);
  and AND2_3708(WX10667,WX10869,WX11348);
  and AND2_3709(WX10668,WX11496,WX10669);
  and AND2_3710(WX10673,WX10684,WX11347);
  and AND2_3711(WX10674,WX10680,WX10675);
  and AND2_3712(WX10677,CRC_OUT_1_10,WX11348);
  and AND2_3713(WX10678,DATA_0_10,WX10679);
  and AND2_3714(WX10681,WX10871,WX11348);
  and AND2_3715(WX10682,WX11503,WX10683);
  and AND2_3716(WX10687,WX10698,WX11347);
  and AND2_3717(WX10688,WX10694,WX10689);
  and AND2_3718(WX10691,CRC_OUT_1_9,WX11348);
  and AND2_3719(WX10692,DATA_0_9,WX10693);
  and AND2_3720(WX10695,WX10873,WX11348);
  and AND2_3721(WX10696,WX11510,WX10697);
  and AND2_3722(WX10701,WX10712,WX11347);
  and AND2_3723(WX10702,WX10708,WX10703);
  and AND2_3724(WX10705,CRC_OUT_1_8,WX11348);
  and AND2_3725(WX10706,DATA_0_8,WX10707);
  and AND2_3726(WX10709,WX10875,WX11348);
  and AND2_3727(WX10710,WX11517,WX10711);
  and AND2_3728(WX10715,WX10726,WX11347);
  and AND2_3729(WX10716,WX10722,WX10717);
  and AND2_3730(WX10719,CRC_OUT_1_7,WX11348);
  and AND2_3731(WX10720,DATA_0_7,WX10721);
  and AND2_3732(WX10723,WX10877,WX11348);
  and AND2_3733(WX10724,WX11524,WX10725);
  and AND2_3734(WX10729,WX10740,WX11347);
  and AND2_3735(WX10730,WX10736,WX10731);
  and AND2_3736(WX10733,CRC_OUT_1_6,WX11348);
  and AND2_3737(WX10734,DATA_0_6,WX10735);
  and AND2_3738(WX10737,WX10879,WX11348);
  and AND2_3739(WX10738,WX11531,WX10739);
  and AND2_3740(WX10743,WX10754,WX11347);
  and AND2_3741(WX10744,WX10750,WX10745);
  and AND2_3742(WX10747,CRC_OUT_1_5,WX11348);
  and AND2_3743(WX10748,DATA_0_5,WX10749);
  and AND2_3744(WX10751,WX10881,WX11348);
  and AND2_3745(WX10752,WX11538,WX10753);
  and AND2_3746(WX10757,WX10768,WX11347);
  and AND2_3747(WX10758,WX10764,WX10759);
  and AND2_3748(WX10761,CRC_OUT_1_4,WX11348);
  and AND2_3749(WX10762,DATA_0_4,WX10763);
  and AND2_3750(WX10765,WX10883,WX11348);
  and AND2_3751(WX10766,WX11545,WX10767);
  and AND2_3752(WX10771,WX10782,WX11347);
  and AND2_3753(WX10772,WX10778,WX10773);
  and AND2_3754(WX10775,CRC_OUT_1_3,WX11348);
  and AND2_3755(WX10776,DATA_0_3,WX10777);
  and AND2_3756(WX10779,WX10885,WX11348);
  and AND2_3757(WX10780,WX11552,WX10781);
  and AND2_3758(WX10785,WX10796,WX11347);
  and AND2_3759(WX10786,WX10792,WX10787);
  and AND2_3760(WX10789,CRC_OUT_1_2,WX11348);
  and AND2_3761(WX10790,DATA_0_2,WX10791);
  and AND2_3762(WX10793,WX10887,WX11348);
  and AND2_3763(WX10794,WX11559,WX10795);
  and AND2_3764(WX10799,WX10810,WX11347);
  and AND2_3765(WX10800,WX10806,WX10801);
  and AND2_3766(WX10803,CRC_OUT_1_1,WX11348);
  and AND2_3767(WX10804,DATA_0_1,WX10805);
  and AND2_3768(WX10807,WX10889,WX11348);
  and AND2_3769(WX10808,WX11566,WX10809);
  and AND2_3770(WX10813,WX10824,WX11347);
  and AND2_3771(WX10814,WX10820,WX10815);
  and AND2_3772(WX10817,CRC_OUT_1_0,WX11348);
  and AND2_3773(WX10818,DATA_0_0,WX10819);
  and AND2_3774(WX10821,WX10891,WX11348);
  and AND2_3775(WX10822,WX11573,WX10823);
  and AND2_3776(WX10828,WX10831,RESET);
  and AND2_3777(WX10830,WX10833,RESET);
  and AND2_3778(WX10832,WX10835,RESET);
  and AND2_3779(WX10834,WX10837,RESET);
  and AND2_3780(WX10836,WX10839,RESET);
  and AND2_3781(WX10838,WX10841,RESET);
  and AND2_3782(WX10840,WX10843,RESET);
  and AND2_3783(WX10842,WX10845,RESET);
  and AND2_3784(WX10844,WX10847,RESET);
  and AND2_3785(WX10846,WX10849,RESET);
  and AND2_3786(WX10848,WX10851,RESET);
  and AND2_3787(WX10850,WX10853,RESET);
  and AND2_3788(WX10852,WX10855,RESET);
  and AND2_3789(WX10854,WX10857,RESET);
  and AND2_3790(WX10856,WX10859,RESET);
  and AND2_3791(WX10858,WX10861,RESET);
  and AND2_3792(WX10860,WX10863,RESET);
  and AND2_3793(WX10862,WX10865,RESET);
  and AND2_3794(WX10864,WX10867,RESET);
  and AND2_3795(WX10866,WX10869,RESET);
  and AND2_3796(WX10868,WX10871,RESET);
  and AND2_3797(WX10870,WX10873,RESET);
  and AND2_3798(WX10872,WX10875,RESET);
  and AND2_3799(WX10874,WX10877,RESET);
  and AND2_3800(WX10876,WX10879,RESET);
  and AND2_3801(WX10878,WX10881,RESET);
  and AND2_3802(WX10880,WX10883,RESET);
  and AND2_3803(WX10882,WX10885,RESET);
  and AND2_3804(WX10884,WX10887,RESET);
  and AND2_3805(WX10886,WX10889,RESET);
  and AND2_3806(WX10888,WX10891,RESET);
  and AND2_3807(WX10890,WX10827,RESET);
  and AND2_3808(WX10988,WX10392,RESET);
  and AND2_3809(WX10990,WX10406,RESET);
  and AND2_3810(WX10992,WX10420,RESET);
  and AND2_3811(WX10994,WX10434,RESET);
  and AND2_3812(WX10996,WX10448,RESET);
  and AND2_3813(WX10998,WX10462,RESET);
  and AND2_3814(WX11000,WX10476,RESET);
  and AND2_3815(WX11002,WX10490,RESET);
  and AND2_3816(WX11004,WX10504,RESET);
  and AND2_3817(WX11006,WX10518,RESET);
  and AND2_3818(WX11008,WX10532,RESET);
  and AND2_3819(WX11010,WX10546,RESET);
  and AND2_3820(WX11012,WX10560,RESET);
  and AND2_3821(WX11014,WX10574,RESET);
  and AND2_3822(WX11016,WX10588,RESET);
  and AND2_3823(WX11018,WX10602,RESET);
  and AND2_3824(WX11020,WX10616,RESET);
  and AND2_3825(WX11022,WX10630,RESET);
  and AND2_3826(WX11024,WX10644,RESET);
  and AND2_3827(WX11026,WX10658,RESET);
  and AND2_3828(WX11028,WX10672,RESET);
  and AND2_3829(WX11030,WX10686,RESET);
  and AND2_3830(WX11032,WX10700,RESET);
  and AND2_3831(WX11034,WX10714,RESET);
  and AND2_3832(WX11036,WX10728,RESET);
  and AND2_3833(WX11038,WX10742,RESET);
  and AND2_3834(WX11040,WX10756,RESET);
  and AND2_3835(WX11042,WX10770,RESET);
  and AND2_3836(WX11044,WX10784,RESET);
  and AND2_3837(WX11046,WX10798,RESET);
  and AND2_3838(WX11048,WX10812,RESET);
  and AND2_3839(WX11050,WX10826,RESET);
  and AND2_3840(WX11052,WX10989,RESET);
  and AND2_3841(WX11054,WX10991,RESET);
  and AND2_3842(WX11056,WX10993,RESET);
  and AND2_3843(WX11058,WX10995,RESET);
  and AND2_3844(WX11060,WX10997,RESET);
  and AND2_3845(WX11062,WX10999,RESET);
  and AND2_3846(WX11064,WX11001,RESET);
  and AND2_3847(WX11066,WX11003,RESET);
  and AND2_3848(WX11068,WX11005,RESET);
  and AND2_3849(WX11070,WX11007,RESET);
  and AND2_3850(WX11072,WX11009,RESET);
  and AND2_3851(WX11074,WX11011,RESET);
  and AND2_3852(WX11076,WX11013,RESET);
  and AND2_3853(WX11078,WX11015,RESET);
  and AND2_3854(WX11080,WX11017,RESET);
  and AND2_3855(WX11082,WX11019,RESET);
  and AND2_3856(WX11084,WX11021,RESET);
  and AND2_3857(WX11086,WX11023,RESET);
  and AND2_3858(WX11088,WX11025,RESET);
  and AND2_3859(WX11090,WX11027,RESET);
  and AND2_3860(WX11092,WX11029,RESET);
  and AND2_3861(WX11094,WX11031,RESET);
  and AND2_3862(WX11096,WX11033,RESET);
  and AND2_3863(WX11098,WX11035,RESET);
  and AND2_3864(WX11100,WX11037,RESET);
  and AND2_3865(WX11102,WX11039,RESET);
  and AND2_3866(WX11104,WX11041,RESET);
  and AND2_3867(WX11106,WX11043,RESET);
  and AND2_3868(WX11108,WX11045,RESET);
  and AND2_3869(WX11110,WX11047,RESET);
  and AND2_3870(WX11112,WX11049,RESET);
  and AND2_3871(WX11114,WX11051,RESET);
  and AND2_3872(WX11116,WX11053,RESET);
  and AND2_3873(WX11118,WX11055,RESET);
  and AND2_3874(WX11120,WX11057,RESET);
  and AND2_3875(WX11122,WX11059,RESET);
  and AND2_3876(WX11124,WX11061,RESET);
  and AND2_3877(WX11126,WX11063,RESET);
  and AND2_3878(WX11128,WX11065,RESET);
  and AND2_3879(WX11130,WX11067,RESET);
  and AND2_3880(WX11132,WX11069,RESET);
  and AND2_3881(WX11134,WX11071,RESET);
  and AND2_3882(WX11136,WX11073,RESET);
  and AND2_3883(WX11138,WX11075,RESET);
  and AND2_3884(WX11140,WX11077,RESET);
  and AND2_3885(WX11142,WX11079,RESET);
  and AND2_3886(WX11144,WX11081,RESET);
  and AND2_3887(WX11146,WX11083,RESET);
  and AND2_3888(WX11148,WX11085,RESET);
  and AND2_3889(WX11150,WX11087,RESET);
  and AND2_3890(WX11152,WX11089,RESET);
  and AND2_3891(WX11154,WX11091,RESET);
  and AND2_3892(WX11156,WX11093,RESET);
  and AND2_3893(WX11158,WX11095,RESET);
  and AND2_3894(WX11160,WX11097,RESET);
  and AND2_3895(WX11162,WX11099,RESET);
  and AND2_3896(WX11164,WX11101,RESET);
  and AND2_3897(WX11166,WX11103,RESET);
  and AND2_3898(WX11168,WX11105,RESET);
  and AND2_3899(WX11170,WX11107,RESET);
  and AND2_3900(WX11172,WX11109,RESET);
  and AND2_3901(WX11174,WX11111,RESET);
  and AND2_3902(WX11176,WX11113,RESET);
  and AND2_3903(WX11178,WX11115,RESET);
  and AND2_3904(WX11180,WX11117,RESET);
  and AND2_3905(WX11182,WX11119,RESET);
  and AND2_3906(WX11184,WX11121,RESET);
  and AND2_3907(WX11186,WX11123,RESET);
  and AND2_3908(WX11188,WX11125,RESET);
  and AND2_3909(WX11190,WX11127,RESET);
  and AND2_3910(WX11192,WX11129,RESET);
  and AND2_3911(WX11194,WX11131,RESET);
  and AND2_3912(WX11196,WX11133,RESET);
  and AND2_3913(WX11198,WX11135,RESET);
  and AND2_3914(WX11200,WX11137,RESET);
  and AND2_3915(WX11202,WX11139,RESET);
  and AND2_3916(WX11204,WX11141,RESET);
  and AND2_3917(WX11206,WX11143,RESET);
  and AND2_3918(WX11208,WX11145,RESET);
  and AND2_3919(WX11210,WX11147,RESET);
  and AND2_3920(WX11212,WX11149,RESET);
  and AND2_3921(WX11214,WX11151,RESET);
  and AND2_3922(WX11216,WX11153,RESET);
  and AND2_3923(WX11218,WX11155,RESET);
  and AND2_3924(WX11220,WX11157,RESET);
  and AND2_3925(WX11222,WX11159,RESET);
  and AND2_3926(WX11224,WX11161,RESET);
  and AND2_3927(WX11226,WX11163,RESET);
  and AND2_3928(WX11228,WX11165,RESET);
  and AND2_3929(WX11230,WX11167,RESET);
  and AND2_3930(WX11232,WX11169,RESET);
  and AND2_3931(WX11234,WX11171,RESET);
  and AND2_3932(WX11236,WX11173,RESET);
  and AND2_3933(WX11238,WX11175,RESET);
  and AND2_3934(WX11240,WX11177,RESET);
  and AND2_3935(WX11242,WX11179,RESET);
  and AND2_3936(WX11351,WX11350,WX11349);
  and AND2_3937(WX11352,WX10924,WX11353);
  and AND2_3938(WX11358,WX11357,WX11349);
  and AND2_3939(WX11359,WX10925,WX11360);
  and AND2_3940(WX11365,WX11364,WX11349);
  and AND2_3941(WX11366,WX10926,WX11367);
  and AND2_3942(WX11372,WX11371,WX11349);
  and AND2_3943(WX11373,WX10927,WX11374);
  and AND2_3944(WX11379,WX11378,WX11349);
  and AND2_3945(WX11380,WX10928,WX11381);
  and AND2_3946(WX11386,WX11385,WX11349);
  and AND2_3947(WX11387,WX10929,WX11388);
  and AND2_3948(WX11393,WX11392,WX11349);
  and AND2_3949(WX11394,WX10930,WX11395);
  and AND2_3950(WX11400,WX11399,WX11349);
  and AND2_3951(WX11401,WX10931,WX11402);
  and AND2_3952(WX11407,WX11406,WX11349);
  and AND2_3953(WX11408,WX10932,WX11409);
  and AND2_3954(WX11414,WX11413,WX11349);
  and AND2_3955(WX11415,WX10933,WX11416);
  and AND2_3956(WX11421,WX11420,WX11349);
  and AND2_3957(WX11422,WX10934,WX11423);
  and AND2_3958(WX11428,WX11427,WX11349);
  and AND2_3959(WX11429,WX10935,WX11430);
  and AND2_3960(WX11435,WX11434,WX11349);
  and AND2_3961(WX11436,WX10936,WX11437);
  and AND2_3962(WX11442,WX11441,WX11349);
  and AND2_3963(WX11443,WX10937,WX11444);
  and AND2_3964(WX11449,WX11448,WX11349);
  and AND2_3965(WX11450,WX10938,WX11451);
  and AND2_3966(WX11456,WX11455,WX11349);
  and AND2_3967(WX11457,WX10939,WX11458);
  and AND2_3968(WX11463,WX11462,WX11349);
  and AND2_3969(WX11464,WX10940,WX11465);
  and AND2_3970(WX11470,WX11469,WX11349);
  and AND2_3971(WX11471,WX10941,WX11472);
  and AND2_3972(WX11477,WX11476,WX11349);
  and AND2_3973(WX11478,WX10942,WX11479);
  and AND2_3974(WX11484,WX11483,WX11349);
  and AND2_3975(WX11485,WX10943,WX11486);
  and AND2_3976(WX11491,WX11490,WX11349);
  and AND2_3977(WX11492,WX10944,WX11493);
  and AND2_3978(WX11498,WX11497,WX11349);
  and AND2_3979(WX11499,WX10945,WX11500);
  and AND2_3980(WX11505,WX11504,WX11349);
  and AND2_3981(WX11506,WX10946,WX11507);
  and AND2_3982(WX11512,WX11511,WX11349);
  and AND2_3983(WX11513,WX10947,WX11514);
  and AND2_3984(WX11519,WX11518,WX11349);
  and AND2_3985(WX11520,WX10948,WX11521);
  and AND2_3986(WX11526,WX11525,WX11349);
  and AND2_3987(WX11527,WX10949,WX11528);
  and AND2_3988(WX11533,WX11532,WX11349);
  and AND2_3989(WX11534,WX10950,WX11535);
  and AND2_3990(WX11540,WX11539,WX11349);
  and AND2_3991(WX11541,WX10951,WX11542);
  and AND2_3992(WX11547,WX11546,WX11349);
  and AND2_3993(WX11548,WX10952,WX11549);
  and AND2_3994(WX11554,WX11553,WX11349);
  and AND2_3995(WX11555,WX10953,WX11556);
  and AND2_3996(WX11561,WX11560,WX11349);
  and AND2_3997(WX11562,WX10954,WX11563);
  and AND2_3998(WX11568,WX11567,WX11349);
  and AND2_3999(WX11569,WX10955,WX11570);
  and AND2_4000(WX11608,WX11578,WX11607);
  and AND2_4001(WX11610,WX11606,WX11607);
  and AND2_4002(WX11612,WX11605,WX11607);
  and AND2_4003(WX11614,WX11604,WX11607);
  and AND2_4004(WX11616,WX11577,WX11607);
  and AND2_4005(WX11618,WX11603,WX11607);
  and AND2_4006(WX11620,WX11602,WX11607);
  and AND2_4007(WX11622,WX11601,WX11607);
  and AND2_4008(WX11624,WX11600,WX11607);
  and AND2_4009(WX11626,WX11599,WX11607);
  and AND2_4010(WX11628,WX11598,WX11607);
  and AND2_4011(WX11630,WX11576,WX11607);
  and AND2_4012(WX11632,WX11597,WX11607);
  and AND2_4013(WX11634,WX11596,WX11607);
  and AND2_4014(WX11636,WX11595,WX11607);
  and AND2_4015(WX11638,WX11594,WX11607);
  and AND2_4016(WX11640,WX11575,WX11607);
  and AND2_4017(WX11642,WX11593,WX11607);
  and AND2_4018(WX11644,WX11592,WX11607);
  and AND2_4019(WX11646,WX11591,WX11607);
  and AND2_4020(WX11648,WX11590,WX11607);
  and AND2_4021(WX11650,WX11589,WX11607);
  and AND2_4022(WX11652,WX11588,WX11607);
  and AND2_4023(WX11654,WX11587,WX11607);
  and AND2_4024(WX11656,WX11586,WX11607);
  and AND2_4025(WX11658,WX11585,WX11607);
  and AND2_4026(WX11660,WX11584,WX11607);
  and AND2_4027(WX11662,WX11583,WX11607);
  and AND2_4028(WX11664,WX11582,WX11607);
  and AND2_4029(WX11666,WX11581,WX11607);
  and AND2_4030(WX11668,WX11580,WX11607);
  and AND2_4031(WX11670,WX11579,WX11607);
  or OR2_0(WX38,WX36,WX35);
  or OR2_1(WX42,WX40,WX39);
  or OR2_2(WX46,WX44,WX43);
  or OR2_3(WX52,WX50,WX49);
  or OR2_4(WX56,WX54,WX53);
  or OR2_5(WX60,WX58,WX57);
  or OR2_6(WX66,WX64,WX63);
  or OR2_7(WX70,WX68,WX67);
  or OR2_8(WX74,WX72,WX71);
  or OR2_9(WX80,WX78,WX77);
  or OR2_10(WX84,WX82,WX81);
  or OR2_11(WX88,WX86,WX85);
  or OR2_12(WX94,WX92,WX91);
  or OR2_13(WX98,WX96,WX95);
  or OR2_14(WX102,WX100,WX99);
  or OR2_15(WX108,WX106,WX105);
  or OR2_16(WX112,WX110,WX109);
  or OR2_17(WX116,WX114,WX113);
  or OR2_18(WX122,WX120,WX119);
  or OR2_19(WX126,WX124,WX123);
  or OR2_20(WX130,WX128,WX127);
  or OR2_21(WX136,WX134,WX133);
  or OR2_22(WX140,WX138,WX137);
  or OR2_23(WX144,WX142,WX141);
  or OR2_24(WX150,WX148,WX147);
  or OR2_25(WX154,WX152,WX151);
  or OR2_26(WX158,WX156,WX155);
  or OR2_27(WX164,WX162,WX161);
  or OR2_28(WX168,WX166,WX165);
  or OR2_29(WX172,WX170,WX169);
  or OR2_30(WX178,WX176,WX175);
  or OR2_31(WX182,WX180,WX179);
  or OR2_32(WX186,WX184,WX183);
  or OR2_33(WX192,WX190,WX189);
  or OR2_34(WX196,WX194,WX193);
  or OR2_35(WX200,WX198,WX197);
  or OR2_36(WX206,WX204,WX203);
  or OR2_37(WX210,WX208,WX207);
  or OR2_38(WX214,WX212,WX211);
  or OR2_39(WX220,WX218,WX217);
  or OR2_40(WX224,WX222,WX221);
  or OR2_41(WX228,WX226,WX225);
  or OR2_42(WX234,WX232,WX231);
  or OR2_43(WX238,WX236,WX235);
  or OR2_44(WX242,WX240,WX239);
  or OR2_45(WX248,WX246,WX245);
  or OR2_46(WX252,WX250,WX249);
  or OR2_47(WX256,WX254,WX253);
  or OR2_48(WX262,WX260,WX259);
  or OR2_49(WX266,WX264,WX263);
  or OR2_50(WX270,WX268,WX267);
  or OR2_51(WX276,WX274,WX273);
  or OR2_52(WX280,WX278,WX277);
  or OR2_53(WX284,WX282,WX281);
  or OR2_54(WX290,WX288,WX287);
  or OR2_55(WX294,WX292,WX291);
  or OR2_56(WX298,WX296,WX295);
  or OR2_57(WX304,WX302,WX301);
  or OR2_58(WX308,WX306,WX305);
  or OR2_59(WX312,WX310,WX309);
  or OR2_60(WX318,WX316,WX315);
  or OR2_61(WX322,WX320,WX319);
  or OR2_62(WX326,WX324,WX323);
  or OR2_63(WX332,WX330,WX329);
  or OR2_64(WX336,WX334,WX333);
  or OR2_65(WX340,WX338,WX337);
  or OR2_66(WX346,WX344,WX343);
  or OR2_67(WX350,WX348,WX347);
  or OR2_68(WX354,WX352,WX351);
  or OR2_69(WX360,WX358,WX357);
  or OR2_70(WX364,WX362,WX361);
  or OR2_71(WX368,WX366,WX365);
  or OR2_72(WX374,WX372,WX371);
  or OR2_73(WX378,WX376,WX375);
  or OR2_74(WX382,WX380,WX379);
  or OR2_75(WX388,WX386,WX385);
  or OR2_76(WX392,WX390,WX389);
  or OR2_77(WX396,WX394,WX393);
  or OR2_78(WX402,WX400,WX399);
  or OR2_79(WX406,WX404,WX403);
  or OR2_80(WX410,WX408,WX407);
  or OR2_81(WX416,WX414,WX413);
  or OR2_82(WX420,WX418,WX417);
  or OR2_83(WX424,WX422,WX421);
  or OR2_84(WX430,WX428,WX427);
  or OR2_85(WX434,WX432,WX431);
  or OR2_86(WX438,WX436,WX435);
  or OR2_87(WX444,WX442,WX441);
  or OR2_88(WX448,WX446,WX445);
  or OR2_89(WX452,WX450,WX449);
  or OR2_90(WX458,WX456,WX455);
  or OR2_91(WX462,WX460,WX459);
  or OR2_92(WX466,WX464,WX463);
  or OR2_93(WX472,WX470,WX469);
  or OR2_94(WX476,WX474,WX473);
  or OR2_95(WX480,WX478,WX477);
  or OR2_96(WX1010,WX1008,WX1007);
  or OR2_97(WX1017,WX1015,WX1014);
  or OR2_98(WX1024,WX1022,WX1021);
  or OR2_99(WX1031,WX1029,WX1028);
  or OR2_100(WX1038,WX1036,WX1035);
  or OR2_101(WX1045,WX1043,WX1042);
  or OR2_102(WX1052,WX1050,WX1049);
  or OR2_103(WX1059,WX1057,WX1056);
  or OR2_104(WX1066,WX1064,WX1063);
  or OR2_105(WX1073,WX1071,WX1070);
  or OR2_106(WX1080,WX1078,WX1077);
  or OR2_107(WX1087,WX1085,WX1084);
  or OR2_108(WX1094,WX1092,WX1091);
  or OR2_109(WX1101,WX1099,WX1098);
  or OR2_110(WX1108,WX1106,WX1105);
  or OR2_111(WX1115,WX1113,WX1112);
  or OR2_112(WX1122,WX1120,WX1119);
  or OR2_113(WX1129,WX1127,WX1126);
  or OR2_114(WX1136,WX1134,WX1133);
  or OR2_115(WX1143,WX1141,WX1140);
  or OR2_116(WX1150,WX1148,WX1147);
  or OR2_117(WX1157,WX1155,WX1154);
  or OR2_118(WX1164,WX1162,WX1161);
  or OR2_119(WX1171,WX1169,WX1168);
  or OR2_120(WX1178,WX1176,WX1175);
  or OR2_121(WX1185,WX1183,WX1182);
  or OR2_122(WX1192,WX1190,WX1189);
  or OR2_123(WX1199,WX1197,WX1196);
  or OR2_124(WX1206,WX1204,WX1203);
  or OR2_125(WX1213,WX1211,WX1210);
  or OR2_126(WX1220,WX1218,WX1217);
  or OR2_127(WX1227,WX1225,WX1224);
  or OR2_128(WX1331,WX1329,WX1328);
  or OR2_129(WX1335,WX1333,WX1332);
  or OR2_130(WX1339,WX1337,WX1336);
  or OR2_131(WX1345,WX1343,WX1342);
  or OR2_132(WX1349,WX1347,WX1346);
  or OR2_133(WX1353,WX1351,WX1350);
  or OR2_134(WX1359,WX1357,WX1356);
  or OR2_135(WX1363,WX1361,WX1360);
  or OR2_136(WX1367,WX1365,WX1364);
  or OR2_137(WX1373,WX1371,WX1370);
  or OR2_138(WX1377,WX1375,WX1374);
  or OR2_139(WX1381,WX1379,WX1378);
  or OR2_140(WX1387,WX1385,WX1384);
  or OR2_141(WX1391,WX1389,WX1388);
  or OR2_142(WX1395,WX1393,WX1392);
  or OR2_143(WX1401,WX1399,WX1398);
  or OR2_144(WX1405,WX1403,WX1402);
  or OR2_145(WX1409,WX1407,WX1406);
  or OR2_146(WX1415,WX1413,WX1412);
  or OR2_147(WX1419,WX1417,WX1416);
  or OR2_148(WX1423,WX1421,WX1420);
  or OR2_149(WX1429,WX1427,WX1426);
  or OR2_150(WX1433,WX1431,WX1430);
  or OR2_151(WX1437,WX1435,WX1434);
  or OR2_152(WX1443,WX1441,WX1440);
  or OR2_153(WX1447,WX1445,WX1444);
  or OR2_154(WX1451,WX1449,WX1448);
  or OR2_155(WX1457,WX1455,WX1454);
  or OR2_156(WX1461,WX1459,WX1458);
  or OR2_157(WX1465,WX1463,WX1462);
  or OR2_158(WX1471,WX1469,WX1468);
  or OR2_159(WX1475,WX1473,WX1472);
  or OR2_160(WX1479,WX1477,WX1476);
  or OR2_161(WX1485,WX1483,WX1482);
  or OR2_162(WX1489,WX1487,WX1486);
  or OR2_163(WX1493,WX1491,WX1490);
  or OR2_164(WX1499,WX1497,WX1496);
  or OR2_165(WX1503,WX1501,WX1500);
  or OR2_166(WX1507,WX1505,WX1504);
  or OR2_167(WX1513,WX1511,WX1510);
  or OR2_168(WX1517,WX1515,WX1514);
  or OR2_169(WX1521,WX1519,WX1518);
  or OR2_170(WX1527,WX1525,WX1524);
  or OR2_171(WX1531,WX1529,WX1528);
  or OR2_172(WX1535,WX1533,WX1532);
  or OR2_173(WX1541,WX1539,WX1538);
  or OR2_174(WX1545,WX1543,WX1542);
  or OR2_175(WX1549,WX1547,WX1546);
  or OR2_176(WX1555,WX1553,WX1552);
  or OR2_177(WX1559,WX1557,WX1556);
  or OR2_178(WX1563,WX1561,WX1560);
  or OR2_179(WX1569,WX1567,WX1566);
  or OR2_180(WX1573,WX1571,WX1570);
  or OR2_181(WX1577,WX1575,WX1574);
  or OR2_182(WX1583,WX1581,WX1580);
  or OR2_183(WX1587,WX1585,WX1584);
  or OR2_184(WX1591,WX1589,WX1588);
  or OR2_185(WX1597,WX1595,WX1594);
  or OR2_186(WX1601,WX1599,WX1598);
  or OR2_187(WX1605,WX1603,WX1602);
  or OR2_188(WX1611,WX1609,WX1608);
  or OR2_189(WX1615,WX1613,WX1612);
  or OR2_190(WX1619,WX1617,WX1616);
  or OR2_191(WX1625,WX1623,WX1622);
  or OR2_192(WX1629,WX1627,WX1626);
  or OR2_193(WX1633,WX1631,WX1630);
  or OR2_194(WX1639,WX1637,WX1636);
  or OR2_195(WX1643,WX1641,WX1640);
  or OR2_196(WX1647,WX1645,WX1644);
  or OR2_197(WX1653,WX1651,WX1650);
  or OR2_198(WX1657,WX1655,WX1654);
  or OR2_199(WX1661,WX1659,WX1658);
  or OR2_200(WX1667,WX1665,WX1664);
  or OR2_201(WX1671,WX1669,WX1668);
  or OR2_202(WX1675,WX1673,WX1672);
  or OR2_203(WX1681,WX1679,WX1678);
  or OR2_204(WX1685,WX1683,WX1682);
  or OR2_205(WX1689,WX1687,WX1686);
  or OR2_206(WX1695,WX1693,WX1692);
  or OR2_207(WX1699,WX1697,WX1696);
  or OR2_208(WX1703,WX1701,WX1700);
  or OR2_209(WX1709,WX1707,WX1706);
  or OR2_210(WX1713,WX1711,WX1710);
  or OR2_211(WX1717,WX1715,WX1714);
  or OR2_212(WX1723,WX1721,WX1720);
  or OR2_213(WX1727,WX1725,WX1724);
  or OR2_214(WX1731,WX1729,WX1728);
  or OR2_215(WX1737,WX1735,WX1734);
  or OR2_216(WX1741,WX1739,WX1738);
  or OR2_217(WX1745,WX1743,WX1742);
  or OR2_218(WX1751,WX1749,WX1748);
  or OR2_219(WX1755,WX1753,WX1752);
  or OR2_220(WX1759,WX1757,WX1756);
  or OR2_221(WX1765,WX1763,WX1762);
  or OR2_222(WX1769,WX1767,WX1766);
  or OR2_223(WX1773,WX1771,WX1770);
  or OR2_224(WX2303,WX2301,WX2300);
  or OR2_225(WX2310,WX2308,WX2307);
  or OR2_226(WX2317,WX2315,WX2314);
  or OR2_227(WX2324,WX2322,WX2321);
  or OR2_228(WX2331,WX2329,WX2328);
  or OR2_229(WX2338,WX2336,WX2335);
  or OR2_230(WX2345,WX2343,WX2342);
  or OR2_231(WX2352,WX2350,WX2349);
  or OR2_232(WX2359,WX2357,WX2356);
  or OR2_233(WX2366,WX2364,WX2363);
  or OR2_234(WX2373,WX2371,WX2370);
  or OR2_235(WX2380,WX2378,WX2377);
  or OR2_236(WX2387,WX2385,WX2384);
  or OR2_237(WX2394,WX2392,WX2391);
  or OR2_238(WX2401,WX2399,WX2398);
  or OR2_239(WX2408,WX2406,WX2405);
  or OR2_240(WX2415,WX2413,WX2412);
  or OR2_241(WX2422,WX2420,WX2419);
  or OR2_242(WX2429,WX2427,WX2426);
  or OR2_243(WX2436,WX2434,WX2433);
  or OR2_244(WX2443,WX2441,WX2440);
  or OR2_245(WX2450,WX2448,WX2447);
  or OR2_246(WX2457,WX2455,WX2454);
  or OR2_247(WX2464,WX2462,WX2461);
  or OR2_248(WX2471,WX2469,WX2468);
  or OR2_249(WX2478,WX2476,WX2475);
  or OR2_250(WX2485,WX2483,WX2482);
  or OR2_251(WX2492,WX2490,WX2489);
  or OR2_252(WX2499,WX2497,WX2496);
  or OR2_253(WX2506,WX2504,WX2503);
  or OR2_254(WX2513,WX2511,WX2510);
  or OR2_255(WX2520,WX2518,WX2517);
  or OR2_256(WX2624,WX2622,WX2621);
  or OR2_257(WX2628,WX2626,WX2625);
  or OR2_258(WX2632,WX2630,WX2629);
  or OR2_259(WX2638,WX2636,WX2635);
  or OR2_260(WX2642,WX2640,WX2639);
  or OR2_261(WX2646,WX2644,WX2643);
  or OR2_262(WX2652,WX2650,WX2649);
  or OR2_263(WX2656,WX2654,WX2653);
  or OR2_264(WX2660,WX2658,WX2657);
  or OR2_265(WX2666,WX2664,WX2663);
  or OR2_266(WX2670,WX2668,WX2667);
  or OR2_267(WX2674,WX2672,WX2671);
  or OR2_268(WX2680,WX2678,WX2677);
  or OR2_269(WX2684,WX2682,WX2681);
  or OR2_270(WX2688,WX2686,WX2685);
  or OR2_271(WX2694,WX2692,WX2691);
  or OR2_272(WX2698,WX2696,WX2695);
  or OR2_273(WX2702,WX2700,WX2699);
  or OR2_274(WX2708,WX2706,WX2705);
  or OR2_275(WX2712,WX2710,WX2709);
  or OR2_276(WX2716,WX2714,WX2713);
  or OR2_277(WX2722,WX2720,WX2719);
  or OR2_278(WX2726,WX2724,WX2723);
  or OR2_279(WX2730,WX2728,WX2727);
  or OR2_280(WX2736,WX2734,WX2733);
  or OR2_281(WX2740,WX2738,WX2737);
  or OR2_282(WX2744,WX2742,WX2741);
  or OR2_283(WX2750,WX2748,WX2747);
  or OR2_284(WX2754,WX2752,WX2751);
  or OR2_285(WX2758,WX2756,WX2755);
  or OR2_286(WX2764,WX2762,WX2761);
  or OR2_287(WX2768,WX2766,WX2765);
  or OR2_288(WX2772,WX2770,WX2769);
  or OR2_289(WX2778,WX2776,WX2775);
  or OR2_290(WX2782,WX2780,WX2779);
  or OR2_291(WX2786,WX2784,WX2783);
  or OR2_292(WX2792,WX2790,WX2789);
  or OR2_293(WX2796,WX2794,WX2793);
  or OR2_294(WX2800,WX2798,WX2797);
  or OR2_295(WX2806,WX2804,WX2803);
  or OR2_296(WX2810,WX2808,WX2807);
  or OR2_297(WX2814,WX2812,WX2811);
  or OR2_298(WX2820,WX2818,WX2817);
  or OR2_299(WX2824,WX2822,WX2821);
  or OR2_300(WX2828,WX2826,WX2825);
  or OR2_301(WX2834,WX2832,WX2831);
  or OR2_302(WX2838,WX2836,WX2835);
  or OR2_303(WX2842,WX2840,WX2839);
  or OR2_304(WX2848,WX2846,WX2845);
  or OR2_305(WX2852,WX2850,WX2849);
  or OR2_306(WX2856,WX2854,WX2853);
  or OR2_307(WX2862,WX2860,WX2859);
  or OR2_308(WX2866,WX2864,WX2863);
  or OR2_309(WX2870,WX2868,WX2867);
  or OR2_310(WX2876,WX2874,WX2873);
  or OR2_311(WX2880,WX2878,WX2877);
  or OR2_312(WX2884,WX2882,WX2881);
  or OR2_313(WX2890,WX2888,WX2887);
  or OR2_314(WX2894,WX2892,WX2891);
  or OR2_315(WX2898,WX2896,WX2895);
  or OR2_316(WX2904,WX2902,WX2901);
  or OR2_317(WX2908,WX2906,WX2905);
  or OR2_318(WX2912,WX2910,WX2909);
  or OR2_319(WX2918,WX2916,WX2915);
  or OR2_320(WX2922,WX2920,WX2919);
  or OR2_321(WX2926,WX2924,WX2923);
  or OR2_322(WX2932,WX2930,WX2929);
  or OR2_323(WX2936,WX2934,WX2933);
  or OR2_324(WX2940,WX2938,WX2937);
  or OR2_325(WX2946,WX2944,WX2943);
  or OR2_326(WX2950,WX2948,WX2947);
  or OR2_327(WX2954,WX2952,WX2951);
  or OR2_328(WX2960,WX2958,WX2957);
  or OR2_329(WX2964,WX2962,WX2961);
  or OR2_330(WX2968,WX2966,WX2965);
  or OR2_331(WX2974,WX2972,WX2971);
  or OR2_332(WX2978,WX2976,WX2975);
  or OR2_333(WX2982,WX2980,WX2979);
  or OR2_334(WX2988,WX2986,WX2985);
  or OR2_335(WX2992,WX2990,WX2989);
  or OR2_336(WX2996,WX2994,WX2993);
  or OR2_337(WX3002,WX3000,WX2999);
  or OR2_338(WX3006,WX3004,WX3003);
  or OR2_339(WX3010,WX3008,WX3007);
  or OR2_340(WX3016,WX3014,WX3013);
  or OR2_341(WX3020,WX3018,WX3017);
  or OR2_342(WX3024,WX3022,WX3021);
  or OR2_343(WX3030,WX3028,WX3027);
  or OR2_344(WX3034,WX3032,WX3031);
  or OR2_345(WX3038,WX3036,WX3035);
  or OR2_346(WX3044,WX3042,WX3041);
  or OR2_347(WX3048,WX3046,WX3045);
  or OR2_348(WX3052,WX3050,WX3049);
  or OR2_349(WX3058,WX3056,WX3055);
  or OR2_350(WX3062,WX3060,WX3059);
  or OR2_351(WX3066,WX3064,WX3063);
  or OR2_352(WX3596,WX3594,WX3593);
  or OR2_353(WX3603,WX3601,WX3600);
  or OR2_354(WX3610,WX3608,WX3607);
  or OR2_355(WX3617,WX3615,WX3614);
  or OR2_356(WX3624,WX3622,WX3621);
  or OR2_357(WX3631,WX3629,WX3628);
  or OR2_358(WX3638,WX3636,WX3635);
  or OR2_359(WX3645,WX3643,WX3642);
  or OR2_360(WX3652,WX3650,WX3649);
  or OR2_361(WX3659,WX3657,WX3656);
  or OR2_362(WX3666,WX3664,WX3663);
  or OR2_363(WX3673,WX3671,WX3670);
  or OR2_364(WX3680,WX3678,WX3677);
  or OR2_365(WX3687,WX3685,WX3684);
  or OR2_366(WX3694,WX3692,WX3691);
  or OR2_367(WX3701,WX3699,WX3698);
  or OR2_368(WX3708,WX3706,WX3705);
  or OR2_369(WX3715,WX3713,WX3712);
  or OR2_370(WX3722,WX3720,WX3719);
  or OR2_371(WX3729,WX3727,WX3726);
  or OR2_372(WX3736,WX3734,WX3733);
  or OR2_373(WX3743,WX3741,WX3740);
  or OR2_374(WX3750,WX3748,WX3747);
  or OR2_375(WX3757,WX3755,WX3754);
  or OR2_376(WX3764,WX3762,WX3761);
  or OR2_377(WX3771,WX3769,WX3768);
  or OR2_378(WX3778,WX3776,WX3775);
  or OR2_379(WX3785,WX3783,WX3782);
  or OR2_380(WX3792,WX3790,WX3789);
  or OR2_381(WX3799,WX3797,WX3796);
  or OR2_382(WX3806,WX3804,WX3803);
  or OR2_383(WX3813,WX3811,WX3810);
  or OR2_384(WX3917,WX3915,WX3914);
  or OR2_385(WX3921,WX3919,WX3918);
  or OR2_386(WX3925,WX3923,WX3922);
  or OR2_387(WX3931,WX3929,WX3928);
  or OR2_388(WX3935,WX3933,WX3932);
  or OR2_389(WX3939,WX3937,WX3936);
  or OR2_390(WX3945,WX3943,WX3942);
  or OR2_391(WX3949,WX3947,WX3946);
  or OR2_392(WX3953,WX3951,WX3950);
  or OR2_393(WX3959,WX3957,WX3956);
  or OR2_394(WX3963,WX3961,WX3960);
  or OR2_395(WX3967,WX3965,WX3964);
  or OR2_396(WX3973,WX3971,WX3970);
  or OR2_397(WX3977,WX3975,WX3974);
  or OR2_398(WX3981,WX3979,WX3978);
  or OR2_399(WX3987,WX3985,WX3984);
  or OR2_400(WX3991,WX3989,WX3988);
  or OR2_401(WX3995,WX3993,WX3992);
  or OR2_402(WX4001,WX3999,WX3998);
  or OR2_403(WX4005,WX4003,WX4002);
  or OR2_404(WX4009,WX4007,WX4006);
  or OR2_405(WX4015,WX4013,WX4012);
  or OR2_406(WX4019,WX4017,WX4016);
  or OR2_407(WX4023,WX4021,WX4020);
  or OR2_408(WX4029,WX4027,WX4026);
  or OR2_409(WX4033,WX4031,WX4030);
  or OR2_410(WX4037,WX4035,WX4034);
  or OR2_411(WX4043,WX4041,WX4040);
  or OR2_412(WX4047,WX4045,WX4044);
  or OR2_413(WX4051,WX4049,WX4048);
  or OR2_414(WX4057,WX4055,WX4054);
  or OR2_415(WX4061,WX4059,WX4058);
  or OR2_416(WX4065,WX4063,WX4062);
  or OR2_417(WX4071,WX4069,WX4068);
  or OR2_418(WX4075,WX4073,WX4072);
  or OR2_419(WX4079,WX4077,WX4076);
  or OR2_420(WX4085,WX4083,WX4082);
  or OR2_421(WX4089,WX4087,WX4086);
  or OR2_422(WX4093,WX4091,WX4090);
  or OR2_423(WX4099,WX4097,WX4096);
  or OR2_424(WX4103,WX4101,WX4100);
  or OR2_425(WX4107,WX4105,WX4104);
  or OR2_426(WX4113,WX4111,WX4110);
  or OR2_427(WX4117,WX4115,WX4114);
  or OR2_428(WX4121,WX4119,WX4118);
  or OR2_429(WX4127,WX4125,WX4124);
  or OR2_430(WX4131,WX4129,WX4128);
  or OR2_431(WX4135,WX4133,WX4132);
  or OR2_432(WX4141,WX4139,WX4138);
  or OR2_433(WX4145,WX4143,WX4142);
  or OR2_434(WX4149,WX4147,WX4146);
  or OR2_435(WX4155,WX4153,WX4152);
  or OR2_436(WX4159,WX4157,WX4156);
  or OR2_437(WX4163,WX4161,WX4160);
  or OR2_438(WX4169,WX4167,WX4166);
  or OR2_439(WX4173,WX4171,WX4170);
  or OR2_440(WX4177,WX4175,WX4174);
  or OR2_441(WX4183,WX4181,WX4180);
  or OR2_442(WX4187,WX4185,WX4184);
  or OR2_443(WX4191,WX4189,WX4188);
  or OR2_444(WX4197,WX4195,WX4194);
  or OR2_445(WX4201,WX4199,WX4198);
  or OR2_446(WX4205,WX4203,WX4202);
  or OR2_447(WX4211,WX4209,WX4208);
  or OR2_448(WX4215,WX4213,WX4212);
  or OR2_449(WX4219,WX4217,WX4216);
  or OR2_450(WX4225,WX4223,WX4222);
  or OR2_451(WX4229,WX4227,WX4226);
  or OR2_452(WX4233,WX4231,WX4230);
  or OR2_453(WX4239,WX4237,WX4236);
  or OR2_454(WX4243,WX4241,WX4240);
  or OR2_455(WX4247,WX4245,WX4244);
  or OR2_456(WX4253,WX4251,WX4250);
  or OR2_457(WX4257,WX4255,WX4254);
  or OR2_458(WX4261,WX4259,WX4258);
  or OR2_459(WX4267,WX4265,WX4264);
  or OR2_460(WX4271,WX4269,WX4268);
  or OR2_461(WX4275,WX4273,WX4272);
  or OR2_462(WX4281,WX4279,WX4278);
  or OR2_463(WX4285,WX4283,WX4282);
  or OR2_464(WX4289,WX4287,WX4286);
  or OR2_465(WX4295,WX4293,WX4292);
  or OR2_466(WX4299,WX4297,WX4296);
  or OR2_467(WX4303,WX4301,WX4300);
  or OR2_468(WX4309,WX4307,WX4306);
  or OR2_469(WX4313,WX4311,WX4310);
  or OR2_470(WX4317,WX4315,WX4314);
  or OR2_471(WX4323,WX4321,WX4320);
  or OR2_472(WX4327,WX4325,WX4324);
  or OR2_473(WX4331,WX4329,WX4328);
  or OR2_474(WX4337,WX4335,WX4334);
  or OR2_475(WX4341,WX4339,WX4338);
  or OR2_476(WX4345,WX4343,WX4342);
  or OR2_477(WX4351,WX4349,WX4348);
  or OR2_478(WX4355,WX4353,WX4352);
  or OR2_479(WX4359,WX4357,WX4356);
  or OR2_480(WX4889,WX4887,WX4886);
  or OR2_481(WX4896,WX4894,WX4893);
  or OR2_482(WX4903,WX4901,WX4900);
  or OR2_483(WX4910,WX4908,WX4907);
  or OR2_484(WX4917,WX4915,WX4914);
  or OR2_485(WX4924,WX4922,WX4921);
  or OR2_486(WX4931,WX4929,WX4928);
  or OR2_487(WX4938,WX4936,WX4935);
  or OR2_488(WX4945,WX4943,WX4942);
  or OR2_489(WX4952,WX4950,WX4949);
  or OR2_490(WX4959,WX4957,WX4956);
  or OR2_491(WX4966,WX4964,WX4963);
  or OR2_492(WX4973,WX4971,WX4970);
  or OR2_493(WX4980,WX4978,WX4977);
  or OR2_494(WX4987,WX4985,WX4984);
  or OR2_495(WX4994,WX4992,WX4991);
  or OR2_496(WX5001,WX4999,WX4998);
  or OR2_497(WX5008,WX5006,WX5005);
  or OR2_498(WX5015,WX5013,WX5012);
  or OR2_499(WX5022,WX5020,WX5019);
  or OR2_500(WX5029,WX5027,WX5026);
  or OR2_501(WX5036,WX5034,WX5033);
  or OR2_502(WX5043,WX5041,WX5040);
  or OR2_503(WX5050,WX5048,WX5047);
  or OR2_504(WX5057,WX5055,WX5054);
  or OR2_505(WX5064,WX5062,WX5061);
  or OR2_506(WX5071,WX5069,WX5068);
  or OR2_507(WX5078,WX5076,WX5075);
  or OR2_508(WX5085,WX5083,WX5082);
  or OR2_509(WX5092,WX5090,WX5089);
  or OR2_510(WX5099,WX5097,WX5096);
  or OR2_511(WX5106,WX5104,WX5103);
  or OR2_512(WX5210,WX5208,WX5207);
  or OR2_513(WX5214,WX5212,WX5211);
  or OR2_514(WX5218,WX5216,WX5215);
  or OR2_515(WX5224,WX5222,WX5221);
  or OR2_516(WX5228,WX5226,WX5225);
  or OR2_517(WX5232,WX5230,WX5229);
  or OR2_518(WX5238,WX5236,WX5235);
  or OR2_519(WX5242,WX5240,WX5239);
  or OR2_520(WX5246,WX5244,WX5243);
  or OR2_521(WX5252,WX5250,WX5249);
  or OR2_522(WX5256,WX5254,WX5253);
  or OR2_523(WX5260,WX5258,WX5257);
  or OR2_524(WX5266,WX5264,WX5263);
  or OR2_525(WX5270,WX5268,WX5267);
  or OR2_526(WX5274,WX5272,WX5271);
  or OR2_527(WX5280,WX5278,WX5277);
  or OR2_528(WX5284,WX5282,WX5281);
  or OR2_529(WX5288,WX5286,WX5285);
  or OR2_530(WX5294,WX5292,WX5291);
  or OR2_531(WX5298,WX5296,WX5295);
  or OR2_532(WX5302,WX5300,WX5299);
  or OR2_533(WX5308,WX5306,WX5305);
  or OR2_534(WX5312,WX5310,WX5309);
  or OR2_535(WX5316,WX5314,WX5313);
  or OR2_536(WX5322,WX5320,WX5319);
  or OR2_537(WX5326,WX5324,WX5323);
  or OR2_538(WX5330,WX5328,WX5327);
  or OR2_539(WX5336,WX5334,WX5333);
  or OR2_540(WX5340,WX5338,WX5337);
  or OR2_541(WX5344,WX5342,WX5341);
  or OR2_542(WX5350,WX5348,WX5347);
  or OR2_543(WX5354,WX5352,WX5351);
  or OR2_544(WX5358,WX5356,WX5355);
  or OR2_545(WX5364,WX5362,WX5361);
  or OR2_546(WX5368,WX5366,WX5365);
  or OR2_547(WX5372,WX5370,WX5369);
  or OR2_548(WX5378,WX5376,WX5375);
  or OR2_549(WX5382,WX5380,WX5379);
  or OR2_550(WX5386,WX5384,WX5383);
  or OR2_551(WX5392,WX5390,WX5389);
  or OR2_552(WX5396,WX5394,WX5393);
  or OR2_553(WX5400,WX5398,WX5397);
  or OR2_554(WX5406,WX5404,WX5403);
  or OR2_555(WX5410,WX5408,WX5407);
  or OR2_556(WX5414,WX5412,WX5411);
  or OR2_557(WX5420,WX5418,WX5417);
  or OR2_558(WX5424,WX5422,WX5421);
  or OR2_559(WX5428,WX5426,WX5425);
  or OR2_560(WX5434,WX5432,WX5431);
  or OR2_561(WX5438,WX5436,WX5435);
  or OR2_562(WX5442,WX5440,WX5439);
  or OR2_563(WX5448,WX5446,WX5445);
  or OR2_564(WX5452,WX5450,WX5449);
  or OR2_565(WX5456,WX5454,WX5453);
  or OR2_566(WX5462,WX5460,WX5459);
  or OR2_567(WX5466,WX5464,WX5463);
  or OR2_568(WX5470,WX5468,WX5467);
  or OR2_569(WX5476,WX5474,WX5473);
  or OR2_570(WX5480,WX5478,WX5477);
  or OR2_571(WX5484,WX5482,WX5481);
  or OR2_572(WX5490,WX5488,WX5487);
  or OR2_573(WX5494,WX5492,WX5491);
  or OR2_574(WX5498,WX5496,WX5495);
  or OR2_575(WX5504,WX5502,WX5501);
  or OR2_576(WX5508,WX5506,WX5505);
  or OR2_577(WX5512,WX5510,WX5509);
  or OR2_578(WX5518,WX5516,WX5515);
  or OR2_579(WX5522,WX5520,WX5519);
  or OR2_580(WX5526,WX5524,WX5523);
  or OR2_581(WX5532,WX5530,WX5529);
  or OR2_582(WX5536,WX5534,WX5533);
  or OR2_583(WX5540,WX5538,WX5537);
  or OR2_584(WX5546,WX5544,WX5543);
  or OR2_585(WX5550,WX5548,WX5547);
  or OR2_586(WX5554,WX5552,WX5551);
  or OR2_587(WX5560,WX5558,WX5557);
  or OR2_588(WX5564,WX5562,WX5561);
  or OR2_589(WX5568,WX5566,WX5565);
  or OR2_590(WX5574,WX5572,WX5571);
  or OR2_591(WX5578,WX5576,WX5575);
  or OR2_592(WX5582,WX5580,WX5579);
  or OR2_593(WX5588,WX5586,WX5585);
  or OR2_594(WX5592,WX5590,WX5589);
  or OR2_595(WX5596,WX5594,WX5593);
  or OR2_596(WX5602,WX5600,WX5599);
  or OR2_597(WX5606,WX5604,WX5603);
  or OR2_598(WX5610,WX5608,WX5607);
  or OR2_599(WX5616,WX5614,WX5613);
  or OR2_600(WX5620,WX5618,WX5617);
  or OR2_601(WX5624,WX5622,WX5621);
  or OR2_602(WX5630,WX5628,WX5627);
  or OR2_603(WX5634,WX5632,WX5631);
  or OR2_604(WX5638,WX5636,WX5635);
  or OR2_605(WX5644,WX5642,WX5641);
  or OR2_606(WX5648,WX5646,WX5645);
  or OR2_607(WX5652,WX5650,WX5649);
  or OR2_608(WX6182,WX6180,WX6179);
  or OR2_609(WX6189,WX6187,WX6186);
  or OR2_610(WX6196,WX6194,WX6193);
  or OR2_611(WX6203,WX6201,WX6200);
  or OR2_612(WX6210,WX6208,WX6207);
  or OR2_613(WX6217,WX6215,WX6214);
  or OR2_614(WX6224,WX6222,WX6221);
  or OR2_615(WX6231,WX6229,WX6228);
  or OR2_616(WX6238,WX6236,WX6235);
  or OR2_617(WX6245,WX6243,WX6242);
  or OR2_618(WX6252,WX6250,WX6249);
  or OR2_619(WX6259,WX6257,WX6256);
  or OR2_620(WX6266,WX6264,WX6263);
  or OR2_621(WX6273,WX6271,WX6270);
  or OR2_622(WX6280,WX6278,WX6277);
  or OR2_623(WX6287,WX6285,WX6284);
  or OR2_624(WX6294,WX6292,WX6291);
  or OR2_625(WX6301,WX6299,WX6298);
  or OR2_626(WX6308,WX6306,WX6305);
  or OR2_627(WX6315,WX6313,WX6312);
  or OR2_628(WX6322,WX6320,WX6319);
  or OR2_629(WX6329,WX6327,WX6326);
  or OR2_630(WX6336,WX6334,WX6333);
  or OR2_631(WX6343,WX6341,WX6340);
  or OR2_632(WX6350,WX6348,WX6347);
  or OR2_633(WX6357,WX6355,WX6354);
  or OR2_634(WX6364,WX6362,WX6361);
  or OR2_635(WX6371,WX6369,WX6368);
  or OR2_636(WX6378,WX6376,WX6375);
  or OR2_637(WX6385,WX6383,WX6382);
  or OR2_638(WX6392,WX6390,WX6389);
  or OR2_639(WX6399,WX6397,WX6396);
  or OR2_640(WX6503,WX6501,WX6500);
  or OR2_641(WX6507,WX6505,WX6504);
  or OR2_642(WX6511,WX6509,WX6508);
  or OR2_643(WX6517,WX6515,WX6514);
  or OR2_644(WX6521,WX6519,WX6518);
  or OR2_645(WX6525,WX6523,WX6522);
  or OR2_646(WX6531,WX6529,WX6528);
  or OR2_647(WX6535,WX6533,WX6532);
  or OR2_648(WX6539,WX6537,WX6536);
  or OR2_649(WX6545,WX6543,WX6542);
  or OR2_650(WX6549,WX6547,WX6546);
  or OR2_651(WX6553,WX6551,WX6550);
  or OR2_652(WX6559,WX6557,WX6556);
  or OR2_653(WX6563,WX6561,WX6560);
  or OR2_654(WX6567,WX6565,WX6564);
  or OR2_655(WX6573,WX6571,WX6570);
  or OR2_656(WX6577,WX6575,WX6574);
  or OR2_657(WX6581,WX6579,WX6578);
  or OR2_658(WX6587,WX6585,WX6584);
  or OR2_659(WX6591,WX6589,WX6588);
  or OR2_660(WX6595,WX6593,WX6592);
  or OR2_661(WX6601,WX6599,WX6598);
  or OR2_662(WX6605,WX6603,WX6602);
  or OR2_663(WX6609,WX6607,WX6606);
  or OR2_664(WX6615,WX6613,WX6612);
  or OR2_665(WX6619,WX6617,WX6616);
  or OR2_666(WX6623,WX6621,WX6620);
  or OR2_667(WX6629,WX6627,WX6626);
  or OR2_668(WX6633,WX6631,WX6630);
  or OR2_669(WX6637,WX6635,WX6634);
  or OR2_670(WX6643,WX6641,WX6640);
  or OR2_671(WX6647,WX6645,WX6644);
  or OR2_672(WX6651,WX6649,WX6648);
  or OR2_673(WX6657,WX6655,WX6654);
  or OR2_674(WX6661,WX6659,WX6658);
  or OR2_675(WX6665,WX6663,WX6662);
  or OR2_676(WX6671,WX6669,WX6668);
  or OR2_677(WX6675,WX6673,WX6672);
  or OR2_678(WX6679,WX6677,WX6676);
  or OR2_679(WX6685,WX6683,WX6682);
  or OR2_680(WX6689,WX6687,WX6686);
  or OR2_681(WX6693,WX6691,WX6690);
  or OR2_682(WX6699,WX6697,WX6696);
  or OR2_683(WX6703,WX6701,WX6700);
  or OR2_684(WX6707,WX6705,WX6704);
  or OR2_685(WX6713,WX6711,WX6710);
  or OR2_686(WX6717,WX6715,WX6714);
  or OR2_687(WX6721,WX6719,WX6718);
  or OR2_688(WX6727,WX6725,WX6724);
  or OR2_689(WX6731,WX6729,WX6728);
  or OR2_690(WX6735,WX6733,WX6732);
  or OR2_691(WX6741,WX6739,WX6738);
  or OR2_692(WX6745,WX6743,WX6742);
  or OR2_693(WX6749,WX6747,WX6746);
  or OR2_694(WX6755,WX6753,WX6752);
  or OR2_695(WX6759,WX6757,WX6756);
  or OR2_696(WX6763,WX6761,WX6760);
  or OR2_697(WX6769,WX6767,WX6766);
  or OR2_698(WX6773,WX6771,WX6770);
  or OR2_699(WX6777,WX6775,WX6774);
  or OR2_700(WX6783,WX6781,WX6780);
  or OR2_701(WX6787,WX6785,WX6784);
  or OR2_702(WX6791,WX6789,WX6788);
  or OR2_703(WX6797,WX6795,WX6794);
  or OR2_704(WX6801,WX6799,WX6798);
  or OR2_705(WX6805,WX6803,WX6802);
  or OR2_706(WX6811,WX6809,WX6808);
  or OR2_707(WX6815,WX6813,WX6812);
  or OR2_708(WX6819,WX6817,WX6816);
  or OR2_709(WX6825,WX6823,WX6822);
  or OR2_710(WX6829,WX6827,WX6826);
  or OR2_711(WX6833,WX6831,WX6830);
  or OR2_712(WX6839,WX6837,WX6836);
  or OR2_713(WX6843,WX6841,WX6840);
  or OR2_714(WX6847,WX6845,WX6844);
  or OR2_715(WX6853,WX6851,WX6850);
  or OR2_716(WX6857,WX6855,WX6854);
  or OR2_717(WX6861,WX6859,WX6858);
  or OR2_718(WX6867,WX6865,WX6864);
  or OR2_719(WX6871,WX6869,WX6868);
  or OR2_720(WX6875,WX6873,WX6872);
  or OR2_721(WX6881,WX6879,WX6878);
  or OR2_722(WX6885,WX6883,WX6882);
  or OR2_723(WX6889,WX6887,WX6886);
  or OR2_724(WX6895,WX6893,WX6892);
  or OR2_725(WX6899,WX6897,WX6896);
  or OR2_726(WX6903,WX6901,WX6900);
  or OR2_727(WX6909,WX6907,WX6906);
  or OR2_728(WX6913,WX6911,WX6910);
  or OR2_729(WX6917,WX6915,WX6914);
  or OR2_730(WX6923,WX6921,WX6920);
  or OR2_731(WX6927,WX6925,WX6924);
  or OR2_732(WX6931,WX6929,WX6928);
  or OR2_733(WX6937,WX6935,WX6934);
  or OR2_734(WX6941,WX6939,WX6938);
  or OR2_735(WX6945,WX6943,WX6942);
  or OR2_736(WX7475,WX7473,WX7472);
  or OR2_737(WX7482,WX7480,WX7479);
  or OR2_738(WX7489,WX7487,WX7486);
  or OR2_739(WX7496,WX7494,WX7493);
  or OR2_740(WX7503,WX7501,WX7500);
  or OR2_741(WX7510,WX7508,WX7507);
  or OR2_742(WX7517,WX7515,WX7514);
  or OR2_743(WX7524,WX7522,WX7521);
  or OR2_744(WX7531,WX7529,WX7528);
  or OR2_745(WX7538,WX7536,WX7535);
  or OR2_746(WX7545,WX7543,WX7542);
  or OR2_747(WX7552,WX7550,WX7549);
  or OR2_748(WX7559,WX7557,WX7556);
  or OR2_749(WX7566,WX7564,WX7563);
  or OR2_750(WX7573,WX7571,WX7570);
  or OR2_751(WX7580,WX7578,WX7577);
  or OR2_752(WX7587,WX7585,WX7584);
  or OR2_753(WX7594,WX7592,WX7591);
  or OR2_754(WX7601,WX7599,WX7598);
  or OR2_755(WX7608,WX7606,WX7605);
  or OR2_756(WX7615,WX7613,WX7612);
  or OR2_757(WX7622,WX7620,WX7619);
  or OR2_758(WX7629,WX7627,WX7626);
  or OR2_759(WX7636,WX7634,WX7633);
  or OR2_760(WX7643,WX7641,WX7640);
  or OR2_761(WX7650,WX7648,WX7647);
  or OR2_762(WX7657,WX7655,WX7654);
  or OR2_763(WX7664,WX7662,WX7661);
  or OR2_764(WX7671,WX7669,WX7668);
  or OR2_765(WX7678,WX7676,WX7675);
  or OR2_766(WX7685,WX7683,WX7682);
  or OR2_767(WX7692,WX7690,WX7689);
  or OR2_768(WX7796,WX7794,WX7793);
  or OR2_769(WX7800,WX7798,WX7797);
  or OR2_770(WX7804,WX7802,WX7801);
  or OR2_771(WX7810,WX7808,WX7807);
  or OR2_772(WX7814,WX7812,WX7811);
  or OR2_773(WX7818,WX7816,WX7815);
  or OR2_774(WX7824,WX7822,WX7821);
  or OR2_775(WX7828,WX7826,WX7825);
  or OR2_776(WX7832,WX7830,WX7829);
  or OR2_777(WX7838,WX7836,WX7835);
  or OR2_778(WX7842,WX7840,WX7839);
  or OR2_779(WX7846,WX7844,WX7843);
  or OR2_780(WX7852,WX7850,WX7849);
  or OR2_781(WX7856,WX7854,WX7853);
  or OR2_782(WX7860,WX7858,WX7857);
  or OR2_783(WX7866,WX7864,WX7863);
  or OR2_784(WX7870,WX7868,WX7867);
  or OR2_785(WX7874,WX7872,WX7871);
  or OR2_786(WX7880,WX7878,WX7877);
  or OR2_787(WX7884,WX7882,WX7881);
  or OR2_788(WX7888,WX7886,WX7885);
  or OR2_789(WX7894,WX7892,WX7891);
  or OR2_790(WX7898,WX7896,WX7895);
  or OR2_791(WX7902,WX7900,WX7899);
  or OR2_792(WX7908,WX7906,WX7905);
  or OR2_793(WX7912,WX7910,WX7909);
  or OR2_794(WX7916,WX7914,WX7913);
  or OR2_795(WX7922,WX7920,WX7919);
  or OR2_796(WX7926,WX7924,WX7923);
  or OR2_797(WX7930,WX7928,WX7927);
  or OR2_798(WX7936,WX7934,WX7933);
  or OR2_799(WX7940,WX7938,WX7937);
  or OR2_800(WX7944,WX7942,WX7941);
  or OR2_801(WX7950,WX7948,WX7947);
  or OR2_802(WX7954,WX7952,WX7951);
  or OR2_803(WX7958,WX7956,WX7955);
  or OR2_804(WX7964,WX7962,WX7961);
  or OR2_805(WX7968,WX7966,WX7965);
  or OR2_806(WX7972,WX7970,WX7969);
  or OR2_807(WX7978,WX7976,WX7975);
  or OR2_808(WX7982,WX7980,WX7979);
  or OR2_809(WX7986,WX7984,WX7983);
  or OR2_810(WX7992,WX7990,WX7989);
  or OR2_811(WX7996,WX7994,WX7993);
  or OR2_812(WX8000,WX7998,WX7997);
  or OR2_813(WX8006,WX8004,WX8003);
  or OR2_814(WX8010,WX8008,WX8007);
  or OR2_815(WX8014,WX8012,WX8011);
  or OR2_816(WX8020,WX8018,WX8017);
  or OR2_817(WX8024,WX8022,WX8021);
  or OR2_818(WX8028,WX8026,WX8025);
  or OR2_819(WX8034,WX8032,WX8031);
  or OR2_820(WX8038,WX8036,WX8035);
  or OR2_821(WX8042,WX8040,WX8039);
  or OR2_822(WX8048,WX8046,WX8045);
  or OR2_823(WX8052,WX8050,WX8049);
  or OR2_824(WX8056,WX8054,WX8053);
  or OR2_825(WX8062,WX8060,WX8059);
  or OR2_826(WX8066,WX8064,WX8063);
  or OR2_827(WX8070,WX8068,WX8067);
  or OR2_828(WX8076,WX8074,WX8073);
  or OR2_829(WX8080,WX8078,WX8077);
  or OR2_830(WX8084,WX8082,WX8081);
  or OR2_831(WX8090,WX8088,WX8087);
  or OR2_832(WX8094,WX8092,WX8091);
  or OR2_833(WX8098,WX8096,WX8095);
  or OR2_834(WX8104,WX8102,WX8101);
  or OR2_835(WX8108,WX8106,WX8105);
  or OR2_836(WX8112,WX8110,WX8109);
  or OR2_837(WX8118,WX8116,WX8115);
  or OR2_838(WX8122,WX8120,WX8119);
  or OR2_839(WX8126,WX8124,WX8123);
  or OR2_840(WX8132,WX8130,WX8129);
  or OR2_841(WX8136,WX8134,WX8133);
  or OR2_842(WX8140,WX8138,WX8137);
  or OR2_843(WX8146,WX8144,WX8143);
  or OR2_844(WX8150,WX8148,WX8147);
  or OR2_845(WX8154,WX8152,WX8151);
  or OR2_846(WX8160,WX8158,WX8157);
  or OR2_847(WX8164,WX8162,WX8161);
  or OR2_848(WX8168,WX8166,WX8165);
  or OR2_849(WX8174,WX8172,WX8171);
  or OR2_850(WX8178,WX8176,WX8175);
  or OR2_851(WX8182,WX8180,WX8179);
  or OR2_852(WX8188,WX8186,WX8185);
  or OR2_853(WX8192,WX8190,WX8189);
  or OR2_854(WX8196,WX8194,WX8193);
  or OR2_855(WX8202,WX8200,WX8199);
  or OR2_856(WX8206,WX8204,WX8203);
  or OR2_857(WX8210,WX8208,WX8207);
  or OR2_858(WX8216,WX8214,WX8213);
  or OR2_859(WX8220,WX8218,WX8217);
  or OR2_860(WX8224,WX8222,WX8221);
  or OR2_861(WX8230,WX8228,WX8227);
  or OR2_862(WX8234,WX8232,WX8231);
  or OR2_863(WX8238,WX8236,WX8235);
  or OR2_864(WX8768,WX8766,WX8765);
  or OR2_865(WX8775,WX8773,WX8772);
  or OR2_866(WX8782,WX8780,WX8779);
  or OR2_867(WX8789,WX8787,WX8786);
  or OR2_868(WX8796,WX8794,WX8793);
  or OR2_869(WX8803,WX8801,WX8800);
  or OR2_870(WX8810,WX8808,WX8807);
  or OR2_871(WX8817,WX8815,WX8814);
  or OR2_872(WX8824,WX8822,WX8821);
  or OR2_873(WX8831,WX8829,WX8828);
  or OR2_874(WX8838,WX8836,WX8835);
  or OR2_875(WX8845,WX8843,WX8842);
  or OR2_876(WX8852,WX8850,WX8849);
  or OR2_877(WX8859,WX8857,WX8856);
  or OR2_878(WX8866,WX8864,WX8863);
  or OR2_879(WX8873,WX8871,WX8870);
  or OR2_880(WX8880,WX8878,WX8877);
  or OR2_881(WX8887,WX8885,WX8884);
  or OR2_882(WX8894,WX8892,WX8891);
  or OR2_883(WX8901,WX8899,WX8898);
  or OR2_884(WX8908,WX8906,WX8905);
  or OR2_885(WX8915,WX8913,WX8912);
  or OR2_886(WX8922,WX8920,WX8919);
  or OR2_887(WX8929,WX8927,WX8926);
  or OR2_888(WX8936,WX8934,WX8933);
  or OR2_889(WX8943,WX8941,WX8940);
  or OR2_890(WX8950,WX8948,WX8947);
  or OR2_891(WX8957,WX8955,WX8954);
  or OR2_892(WX8964,WX8962,WX8961);
  or OR2_893(WX8971,WX8969,WX8968);
  or OR2_894(WX8978,WX8976,WX8975);
  or OR2_895(WX8985,WX8983,WX8982);
  or OR2_896(WX9089,WX9087,WX9086);
  or OR2_897(WX9093,WX9091,WX9090);
  or OR2_898(WX9097,WX9095,WX9094);
  or OR2_899(WX9103,WX9101,WX9100);
  or OR2_900(WX9107,WX9105,WX9104);
  or OR2_901(WX9111,WX9109,WX9108);
  or OR2_902(WX9117,WX9115,WX9114);
  or OR2_903(WX9121,WX9119,WX9118);
  or OR2_904(WX9125,WX9123,WX9122);
  or OR2_905(WX9131,WX9129,WX9128);
  or OR2_906(WX9135,WX9133,WX9132);
  or OR2_907(WX9139,WX9137,WX9136);
  or OR2_908(WX9145,WX9143,WX9142);
  or OR2_909(WX9149,WX9147,WX9146);
  or OR2_910(WX9153,WX9151,WX9150);
  or OR2_911(WX9159,WX9157,WX9156);
  or OR2_912(WX9163,WX9161,WX9160);
  or OR2_913(WX9167,WX9165,WX9164);
  or OR2_914(WX9173,WX9171,WX9170);
  or OR2_915(WX9177,WX9175,WX9174);
  or OR2_916(WX9181,WX9179,WX9178);
  or OR2_917(WX9187,WX9185,WX9184);
  or OR2_918(WX9191,WX9189,WX9188);
  or OR2_919(WX9195,WX9193,WX9192);
  or OR2_920(WX9201,WX9199,WX9198);
  or OR2_921(WX9205,WX9203,WX9202);
  or OR2_922(WX9209,WX9207,WX9206);
  or OR2_923(WX9215,WX9213,WX9212);
  or OR2_924(WX9219,WX9217,WX9216);
  or OR2_925(WX9223,WX9221,WX9220);
  or OR2_926(WX9229,WX9227,WX9226);
  or OR2_927(WX9233,WX9231,WX9230);
  or OR2_928(WX9237,WX9235,WX9234);
  or OR2_929(WX9243,WX9241,WX9240);
  or OR2_930(WX9247,WX9245,WX9244);
  or OR2_931(WX9251,WX9249,WX9248);
  or OR2_932(WX9257,WX9255,WX9254);
  or OR2_933(WX9261,WX9259,WX9258);
  or OR2_934(WX9265,WX9263,WX9262);
  or OR2_935(WX9271,WX9269,WX9268);
  or OR2_936(WX9275,WX9273,WX9272);
  or OR2_937(WX9279,WX9277,WX9276);
  or OR2_938(WX9285,WX9283,WX9282);
  or OR2_939(WX9289,WX9287,WX9286);
  or OR2_940(WX9293,WX9291,WX9290);
  or OR2_941(WX9299,WX9297,WX9296);
  or OR2_942(WX9303,WX9301,WX9300);
  or OR2_943(WX9307,WX9305,WX9304);
  or OR2_944(WX9313,WX9311,WX9310);
  or OR2_945(WX9317,WX9315,WX9314);
  or OR2_946(WX9321,WX9319,WX9318);
  or OR2_947(WX9327,WX9325,WX9324);
  or OR2_948(WX9331,WX9329,WX9328);
  or OR2_949(WX9335,WX9333,WX9332);
  or OR2_950(WX9341,WX9339,WX9338);
  or OR2_951(WX9345,WX9343,WX9342);
  or OR2_952(WX9349,WX9347,WX9346);
  or OR2_953(WX9355,WX9353,WX9352);
  or OR2_954(WX9359,WX9357,WX9356);
  or OR2_955(WX9363,WX9361,WX9360);
  or OR2_956(WX9369,WX9367,WX9366);
  or OR2_957(WX9373,WX9371,WX9370);
  or OR2_958(WX9377,WX9375,WX9374);
  or OR2_959(WX9383,WX9381,WX9380);
  or OR2_960(WX9387,WX9385,WX9384);
  or OR2_961(WX9391,WX9389,WX9388);
  or OR2_962(WX9397,WX9395,WX9394);
  or OR2_963(WX9401,WX9399,WX9398);
  or OR2_964(WX9405,WX9403,WX9402);
  or OR2_965(WX9411,WX9409,WX9408);
  or OR2_966(WX9415,WX9413,WX9412);
  or OR2_967(WX9419,WX9417,WX9416);
  or OR2_968(WX9425,WX9423,WX9422);
  or OR2_969(WX9429,WX9427,WX9426);
  or OR2_970(WX9433,WX9431,WX9430);
  or OR2_971(WX9439,WX9437,WX9436);
  or OR2_972(WX9443,WX9441,WX9440);
  or OR2_973(WX9447,WX9445,WX9444);
  or OR2_974(WX9453,WX9451,WX9450);
  or OR2_975(WX9457,WX9455,WX9454);
  or OR2_976(WX9461,WX9459,WX9458);
  or OR2_977(WX9467,WX9465,WX9464);
  or OR2_978(WX9471,WX9469,WX9468);
  or OR2_979(WX9475,WX9473,WX9472);
  or OR2_980(WX9481,WX9479,WX9478);
  or OR2_981(WX9485,WX9483,WX9482);
  or OR2_982(WX9489,WX9487,WX9486);
  or OR2_983(WX9495,WX9493,WX9492);
  or OR2_984(WX9499,WX9497,WX9496);
  or OR2_985(WX9503,WX9501,WX9500);
  or OR2_986(WX9509,WX9507,WX9506);
  or OR2_987(WX9513,WX9511,WX9510);
  or OR2_988(WX9517,WX9515,WX9514);
  or OR2_989(WX9523,WX9521,WX9520);
  or OR2_990(WX9527,WX9525,WX9524);
  or OR2_991(WX9531,WX9529,WX9528);
  or OR2_992(WX10061,WX10059,WX10058);
  or OR2_993(WX10068,WX10066,WX10065);
  or OR2_994(WX10075,WX10073,WX10072);
  or OR2_995(WX10082,WX10080,WX10079);
  or OR2_996(WX10089,WX10087,WX10086);
  or OR2_997(WX10096,WX10094,WX10093);
  or OR2_998(WX10103,WX10101,WX10100);
  or OR2_999(WX10110,WX10108,WX10107);
  or OR2_1000(WX10117,WX10115,WX10114);
  or OR2_1001(WX10124,WX10122,WX10121);
  or OR2_1002(WX10131,WX10129,WX10128);
  or OR2_1003(WX10138,WX10136,WX10135);
  or OR2_1004(WX10145,WX10143,WX10142);
  or OR2_1005(WX10152,WX10150,WX10149);
  or OR2_1006(WX10159,WX10157,WX10156);
  or OR2_1007(WX10166,WX10164,WX10163);
  or OR2_1008(WX10173,WX10171,WX10170);
  or OR2_1009(WX10180,WX10178,WX10177);
  or OR2_1010(WX10187,WX10185,WX10184);
  or OR2_1011(WX10194,WX10192,WX10191);
  or OR2_1012(WX10201,WX10199,WX10198);
  or OR2_1013(WX10208,WX10206,WX10205);
  or OR2_1014(WX10215,WX10213,WX10212);
  or OR2_1015(WX10222,WX10220,WX10219);
  or OR2_1016(WX10229,WX10227,WX10226);
  or OR2_1017(WX10236,WX10234,WX10233);
  or OR2_1018(WX10243,WX10241,WX10240);
  or OR2_1019(WX10250,WX10248,WX10247);
  or OR2_1020(WX10257,WX10255,WX10254);
  or OR2_1021(WX10264,WX10262,WX10261);
  or OR2_1022(WX10271,WX10269,WX10268);
  or OR2_1023(WX10278,WX10276,WX10275);
  or OR2_1024(WX10382,WX10380,WX10379);
  or OR2_1025(WX10386,WX10384,WX10383);
  or OR2_1026(WX10390,WX10388,WX10387);
  or OR2_1027(WX10396,WX10394,WX10393);
  or OR2_1028(WX10400,WX10398,WX10397);
  or OR2_1029(WX10404,WX10402,WX10401);
  or OR2_1030(WX10410,WX10408,WX10407);
  or OR2_1031(WX10414,WX10412,WX10411);
  or OR2_1032(WX10418,WX10416,WX10415);
  or OR2_1033(WX10424,WX10422,WX10421);
  or OR2_1034(WX10428,WX10426,WX10425);
  or OR2_1035(WX10432,WX10430,WX10429);
  or OR2_1036(WX10438,WX10436,WX10435);
  or OR2_1037(WX10442,WX10440,WX10439);
  or OR2_1038(WX10446,WX10444,WX10443);
  or OR2_1039(WX10452,WX10450,WX10449);
  or OR2_1040(WX10456,WX10454,WX10453);
  or OR2_1041(WX10460,WX10458,WX10457);
  or OR2_1042(WX10466,WX10464,WX10463);
  or OR2_1043(WX10470,WX10468,WX10467);
  or OR2_1044(WX10474,WX10472,WX10471);
  or OR2_1045(WX10480,WX10478,WX10477);
  or OR2_1046(WX10484,WX10482,WX10481);
  or OR2_1047(WX10488,WX10486,WX10485);
  or OR2_1048(WX10494,WX10492,WX10491);
  or OR2_1049(WX10498,WX10496,WX10495);
  or OR2_1050(WX10502,WX10500,WX10499);
  or OR2_1051(WX10508,WX10506,WX10505);
  or OR2_1052(WX10512,WX10510,WX10509);
  or OR2_1053(WX10516,WX10514,WX10513);
  or OR2_1054(WX10522,WX10520,WX10519);
  or OR2_1055(WX10526,WX10524,WX10523);
  or OR2_1056(WX10530,WX10528,WX10527);
  or OR2_1057(WX10536,WX10534,WX10533);
  or OR2_1058(WX10540,WX10538,WX10537);
  or OR2_1059(WX10544,WX10542,WX10541);
  or OR2_1060(WX10550,WX10548,WX10547);
  or OR2_1061(WX10554,WX10552,WX10551);
  or OR2_1062(WX10558,WX10556,WX10555);
  or OR2_1063(WX10564,WX10562,WX10561);
  or OR2_1064(WX10568,WX10566,WX10565);
  or OR2_1065(WX10572,WX10570,WX10569);
  or OR2_1066(WX10578,WX10576,WX10575);
  or OR2_1067(WX10582,WX10580,WX10579);
  or OR2_1068(WX10586,WX10584,WX10583);
  or OR2_1069(WX10592,WX10590,WX10589);
  or OR2_1070(WX10596,WX10594,WX10593);
  or OR2_1071(WX10600,WX10598,WX10597);
  or OR2_1072(WX10606,WX10604,WX10603);
  or OR2_1073(WX10610,WX10608,WX10607);
  or OR2_1074(WX10614,WX10612,WX10611);
  or OR2_1075(WX10620,WX10618,WX10617);
  or OR2_1076(WX10624,WX10622,WX10621);
  or OR2_1077(WX10628,WX10626,WX10625);
  or OR2_1078(WX10634,WX10632,WX10631);
  or OR2_1079(WX10638,WX10636,WX10635);
  or OR2_1080(WX10642,WX10640,WX10639);
  or OR2_1081(WX10648,WX10646,WX10645);
  or OR2_1082(WX10652,WX10650,WX10649);
  or OR2_1083(WX10656,WX10654,WX10653);
  or OR2_1084(WX10662,WX10660,WX10659);
  or OR2_1085(WX10666,WX10664,WX10663);
  or OR2_1086(WX10670,WX10668,WX10667);
  or OR2_1087(WX10676,WX10674,WX10673);
  or OR2_1088(WX10680,WX10678,WX10677);
  or OR2_1089(WX10684,WX10682,WX10681);
  or OR2_1090(WX10690,WX10688,WX10687);
  or OR2_1091(WX10694,WX10692,WX10691);
  or OR2_1092(WX10698,WX10696,WX10695);
  or OR2_1093(WX10704,WX10702,WX10701);
  or OR2_1094(WX10708,WX10706,WX10705);
  or OR2_1095(WX10712,WX10710,WX10709);
  or OR2_1096(WX10718,WX10716,WX10715);
  or OR2_1097(WX10722,WX10720,WX10719);
  or OR2_1098(WX10726,WX10724,WX10723);
  or OR2_1099(WX10732,WX10730,WX10729);
  or OR2_1100(WX10736,WX10734,WX10733);
  or OR2_1101(WX10740,WX10738,WX10737);
  or OR2_1102(WX10746,WX10744,WX10743);
  or OR2_1103(WX10750,WX10748,WX10747);
  or OR2_1104(WX10754,WX10752,WX10751);
  or OR2_1105(WX10760,WX10758,WX10757);
  or OR2_1106(WX10764,WX10762,WX10761);
  or OR2_1107(WX10768,WX10766,WX10765);
  or OR2_1108(WX10774,WX10772,WX10771);
  or OR2_1109(WX10778,WX10776,WX10775);
  or OR2_1110(WX10782,WX10780,WX10779);
  or OR2_1111(WX10788,WX10786,WX10785);
  or OR2_1112(WX10792,WX10790,WX10789);
  or OR2_1113(WX10796,WX10794,WX10793);
  or OR2_1114(WX10802,WX10800,WX10799);
  or OR2_1115(WX10806,WX10804,WX10803);
  or OR2_1116(WX10810,WX10808,WX10807);
  or OR2_1117(WX10816,WX10814,WX10813);
  or OR2_1118(WX10820,WX10818,WX10817);
  or OR2_1119(WX10824,WX10822,WX10821);
  or OR2_1120(WX11354,WX11352,WX11351);
  or OR2_1121(WX11361,WX11359,WX11358);
  or OR2_1122(WX11368,WX11366,WX11365);
  or OR2_1123(WX11375,WX11373,WX11372);
  or OR2_1124(WX11382,WX11380,WX11379);
  or OR2_1125(WX11389,WX11387,WX11386);
  or OR2_1126(WX11396,WX11394,WX11393);
  or OR2_1127(WX11403,WX11401,WX11400);
  or OR2_1128(WX11410,WX11408,WX11407);
  or OR2_1129(WX11417,WX11415,WX11414);
  or OR2_1130(WX11424,WX11422,WX11421);
  or OR2_1131(WX11431,WX11429,WX11428);
  or OR2_1132(WX11438,WX11436,WX11435);
  or OR2_1133(WX11445,WX11443,WX11442);
  or OR2_1134(WX11452,WX11450,WX11449);
  or OR2_1135(WX11459,WX11457,WX11456);
  or OR2_1136(WX11466,WX11464,WX11463);
  or OR2_1137(WX11473,WX11471,WX11470);
  or OR2_1138(WX11480,WX11478,WX11477);
  or OR2_1139(WX11487,WX11485,WX11484);
  or OR2_1140(WX11494,WX11492,WX11491);
  or OR2_1141(WX11501,WX11499,WX11498);
  or OR2_1142(WX11508,WX11506,WX11505);
  or OR2_1143(WX11515,WX11513,WX11512);
  or OR2_1144(WX11522,WX11520,WX11519);
  or OR2_1145(WX11529,WX11527,WX11526);
  or OR2_1146(WX11536,WX11534,WX11533);
  or OR2_1147(WX11543,WX11541,WX11540);
  or OR2_1148(WX11550,WX11548,WX11547);
  or OR2_1149(WX11557,WX11555,WX11554);
  or OR2_1150(WX11564,WX11562,WX11561);
  or OR2_1151(WX11571,WX11569,WX11568);
  nand NAND2_0(II1988,WX1001,WX645);
  nand NAND2_1(II1989,WX1001,II1988);
  nand NAND2_2(II1990,WX645,II1988);
  nand NAND2_3(II1987,II1989,II1990);
  nand NAND2_4(II1995,WX709,II1987);
  nand NAND2_5(II1996,WX709,II1995);
  nand NAND2_6(II1997,II1987,II1995);
  nand NAND2_7(II1986,II1996,II1997);
  nand NAND2_8(II2003,WX773,WX837);
  nand NAND2_9(II2004,WX773,II2003);
  nand NAND2_10(II2005,WX837,II2003);
  nand NAND2_11(II2002,II2004,II2005);
  nand NAND2_12(II2010,II1986,II2002);
  nand NAND2_13(II2011,II1986,II2010);
  nand NAND2_14(II2012,II2002,II2010);
  nand NAND2_15(WX900,II2011,II2012);
  nand NAND2_16(II2019,WX1001,WX647);
  nand NAND2_17(II2020,WX1001,II2019);
  nand NAND2_18(II2021,WX647,II2019);
  nand NAND2_19(II2018,II2020,II2021);
  nand NAND2_20(II2026,WX711,II2018);
  nand NAND2_21(II2027,WX711,II2026);
  nand NAND2_22(II2028,II2018,II2026);
  nand NAND2_23(II2017,II2027,II2028);
  nand NAND2_24(II2034,WX775,WX839);
  nand NAND2_25(II2035,WX775,II2034);
  nand NAND2_26(II2036,WX839,II2034);
  nand NAND2_27(II2033,II2035,II2036);
  nand NAND2_28(II2041,II2017,II2033);
  nand NAND2_29(II2042,II2017,II2041);
  nand NAND2_30(II2043,II2033,II2041);
  nand NAND2_31(WX901,II2042,II2043);
  nand NAND2_32(II2050,WX1001,WX649);
  nand NAND2_33(II2051,WX1001,II2050);
  nand NAND2_34(II2052,WX649,II2050);
  nand NAND2_35(II2049,II2051,II2052);
  nand NAND2_36(II2057,WX713,II2049);
  nand NAND2_37(II2058,WX713,II2057);
  nand NAND2_38(II2059,II2049,II2057);
  nand NAND2_39(II2048,II2058,II2059);
  nand NAND2_40(II2065,WX777,WX841);
  nand NAND2_41(II2066,WX777,II2065);
  nand NAND2_42(II2067,WX841,II2065);
  nand NAND2_43(II2064,II2066,II2067);
  nand NAND2_44(II2072,II2048,II2064);
  nand NAND2_45(II2073,II2048,II2072);
  nand NAND2_46(II2074,II2064,II2072);
  nand NAND2_47(WX902,II2073,II2074);
  nand NAND2_48(II2081,WX1001,WX651);
  nand NAND2_49(II2082,WX1001,II2081);
  nand NAND2_50(II2083,WX651,II2081);
  nand NAND2_51(II2080,II2082,II2083);
  nand NAND2_52(II2088,WX715,II2080);
  nand NAND2_53(II2089,WX715,II2088);
  nand NAND2_54(II2090,II2080,II2088);
  nand NAND2_55(II2079,II2089,II2090);
  nand NAND2_56(II2096,WX779,WX843);
  nand NAND2_57(II2097,WX779,II2096);
  nand NAND2_58(II2098,WX843,II2096);
  nand NAND2_59(II2095,II2097,II2098);
  nand NAND2_60(II2103,II2079,II2095);
  nand NAND2_61(II2104,II2079,II2103);
  nand NAND2_62(II2105,II2095,II2103);
  nand NAND2_63(WX903,II2104,II2105);
  nand NAND2_64(II2112,WX1001,WX653);
  nand NAND2_65(II2113,WX1001,II2112);
  nand NAND2_66(II2114,WX653,II2112);
  nand NAND2_67(II2111,II2113,II2114);
  nand NAND2_68(II2119,WX717,II2111);
  nand NAND2_69(II2120,WX717,II2119);
  nand NAND2_70(II2121,II2111,II2119);
  nand NAND2_71(II2110,II2120,II2121);
  nand NAND2_72(II2127,WX781,WX845);
  nand NAND2_73(II2128,WX781,II2127);
  nand NAND2_74(II2129,WX845,II2127);
  nand NAND2_75(II2126,II2128,II2129);
  nand NAND2_76(II2134,II2110,II2126);
  nand NAND2_77(II2135,II2110,II2134);
  nand NAND2_78(II2136,II2126,II2134);
  nand NAND2_79(WX904,II2135,II2136);
  nand NAND2_80(II2143,WX1001,WX655);
  nand NAND2_81(II2144,WX1001,II2143);
  nand NAND2_82(II2145,WX655,II2143);
  nand NAND2_83(II2142,II2144,II2145);
  nand NAND2_84(II2150,WX719,II2142);
  nand NAND2_85(II2151,WX719,II2150);
  nand NAND2_86(II2152,II2142,II2150);
  nand NAND2_87(II2141,II2151,II2152);
  nand NAND2_88(II2158,WX783,WX847);
  nand NAND2_89(II2159,WX783,II2158);
  nand NAND2_90(II2160,WX847,II2158);
  nand NAND2_91(II2157,II2159,II2160);
  nand NAND2_92(II2165,II2141,II2157);
  nand NAND2_93(II2166,II2141,II2165);
  nand NAND2_94(II2167,II2157,II2165);
  nand NAND2_95(WX905,II2166,II2167);
  nand NAND2_96(II2174,WX1001,WX657);
  nand NAND2_97(II2175,WX1001,II2174);
  nand NAND2_98(II2176,WX657,II2174);
  nand NAND2_99(II2173,II2175,II2176);
  nand NAND2_100(II2181,WX721,II2173);
  nand NAND2_101(II2182,WX721,II2181);
  nand NAND2_102(II2183,II2173,II2181);
  nand NAND2_103(II2172,II2182,II2183);
  nand NAND2_104(II2189,WX785,WX849);
  nand NAND2_105(II2190,WX785,II2189);
  nand NAND2_106(II2191,WX849,II2189);
  nand NAND2_107(II2188,II2190,II2191);
  nand NAND2_108(II2196,II2172,II2188);
  nand NAND2_109(II2197,II2172,II2196);
  nand NAND2_110(II2198,II2188,II2196);
  nand NAND2_111(WX906,II2197,II2198);
  nand NAND2_112(II2205,WX1001,WX659);
  nand NAND2_113(II2206,WX1001,II2205);
  nand NAND2_114(II2207,WX659,II2205);
  nand NAND2_115(II2204,II2206,II2207);
  nand NAND2_116(II2212,WX723,II2204);
  nand NAND2_117(II2213,WX723,II2212);
  nand NAND2_118(II2214,II2204,II2212);
  nand NAND2_119(II2203,II2213,II2214);
  nand NAND2_120(II2220,WX787,WX851);
  nand NAND2_121(II2221,WX787,II2220);
  nand NAND2_122(II2222,WX851,II2220);
  nand NAND2_123(II2219,II2221,II2222);
  nand NAND2_124(II2227,II2203,II2219);
  nand NAND2_125(II2228,II2203,II2227);
  nand NAND2_126(II2229,II2219,II2227);
  nand NAND2_127(WX907,II2228,II2229);
  nand NAND2_128(II2236,WX1001,WX661);
  nand NAND2_129(II2237,WX1001,II2236);
  nand NAND2_130(II2238,WX661,II2236);
  nand NAND2_131(II2235,II2237,II2238);
  nand NAND2_132(II2243,WX725,II2235);
  nand NAND2_133(II2244,WX725,II2243);
  nand NAND2_134(II2245,II2235,II2243);
  nand NAND2_135(II2234,II2244,II2245);
  nand NAND2_136(II2251,WX789,WX853);
  nand NAND2_137(II2252,WX789,II2251);
  nand NAND2_138(II2253,WX853,II2251);
  nand NAND2_139(II2250,II2252,II2253);
  nand NAND2_140(II2258,II2234,II2250);
  nand NAND2_141(II2259,II2234,II2258);
  nand NAND2_142(II2260,II2250,II2258);
  nand NAND2_143(WX908,II2259,II2260);
  nand NAND2_144(II2267,WX1001,WX663);
  nand NAND2_145(II2268,WX1001,II2267);
  nand NAND2_146(II2269,WX663,II2267);
  nand NAND2_147(II2266,II2268,II2269);
  nand NAND2_148(II2274,WX727,II2266);
  nand NAND2_149(II2275,WX727,II2274);
  nand NAND2_150(II2276,II2266,II2274);
  nand NAND2_151(II2265,II2275,II2276);
  nand NAND2_152(II2282,WX791,WX855);
  nand NAND2_153(II2283,WX791,II2282);
  nand NAND2_154(II2284,WX855,II2282);
  nand NAND2_155(II2281,II2283,II2284);
  nand NAND2_156(II2289,II2265,II2281);
  nand NAND2_157(II2290,II2265,II2289);
  nand NAND2_158(II2291,II2281,II2289);
  nand NAND2_159(WX909,II2290,II2291);
  nand NAND2_160(II2298,WX1001,WX665);
  nand NAND2_161(II2299,WX1001,II2298);
  nand NAND2_162(II2300,WX665,II2298);
  nand NAND2_163(II2297,II2299,II2300);
  nand NAND2_164(II2305,WX729,II2297);
  nand NAND2_165(II2306,WX729,II2305);
  nand NAND2_166(II2307,II2297,II2305);
  nand NAND2_167(II2296,II2306,II2307);
  nand NAND2_168(II2313,WX793,WX857);
  nand NAND2_169(II2314,WX793,II2313);
  nand NAND2_170(II2315,WX857,II2313);
  nand NAND2_171(II2312,II2314,II2315);
  nand NAND2_172(II2320,II2296,II2312);
  nand NAND2_173(II2321,II2296,II2320);
  nand NAND2_174(II2322,II2312,II2320);
  nand NAND2_175(WX910,II2321,II2322);
  nand NAND2_176(II2329,WX1001,WX667);
  nand NAND2_177(II2330,WX1001,II2329);
  nand NAND2_178(II2331,WX667,II2329);
  nand NAND2_179(II2328,II2330,II2331);
  nand NAND2_180(II2336,WX731,II2328);
  nand NAND2_181(II2337,WX731,II2336);
  nand NAND2_182(II2338,II2328,II2336);
  nand NAND2_183(II2327,II2337,II2338);
  nand NAND2_184(II2344,WX795,WX859);
  nand NAND2_185(II2345,WX795,II2344);
  nand NAND2_186(II2346,WX859,II2344);
  nand NAND2_187(II2343,II2345,II2346);
  nand NAND2_188(II2351,II2327,II2343);
  nand NAND2_189(II2352,II2327,II2351);
  nand NAND2_190(II2353,II2343,II2351);
  nand NAND2_191(WX911,II2352,II2353);
  nand NAND2_192(II2360,WX1001,WX669);
  nand NAND2_193(II2361,WX1001,II2360);
  nand NAND2_194(II2362,WX669,II2360);
  nand NAND2_195(II2359,II2361,II2362);
  nand NAND2_196(II2367,WX733,II2359);
  nand NAND2_197(II2368,WX733,II2367);
  nand NAND2_198(II2369,II2359,II2367);
  nand NAND2_199(II2358,II2368,II2369);
  nand NAND2_200(II2375,WX797,WX861);
  nand NAND2_201(II2376,WX797,II2375);
  nand NAND2_202(II2377,WX861,II2375);
  nand NAND2_203(II2374,II2376,II2377);
  nand NAND2_204(II2382,II2358,II2374);
  nand NAND2_205(II2383,II2358,II2382);
  nand NAND2_206(II2384,II2374,II2382);
  nand NAND2_207(WX912,II2383,II2384);
  nand NAND2_208(II2391,WX1001,WX671);
  nand NAND2_209(II2392,WX1001,II2391);
  nand NAND2_210(II2393,WX671,II2391);
  nand NAND2_211(II2390,II2392,II2393);
  nand NAND2_212(II2398,WX735,II2390);
  nand NAND2_213(II2399,WX735,II2398);
  nand NAND2_214(II2400,II2390,II2398);
  nand NAND2_215(II2389,II2399,II2400);
  nand NAND2_216(II2406,WX799,WX863);
  nand NAND2_217(II2407,WX799,II2406);
  nand NAND2_218(II2408,WX863,II2406);
  nand NAND2_219(II2405,II2407,II2408);
  nand NAND2_220(II2413,II2389,II2405);
  nand NAND2_221(II2414,II2389,II2413);
  nand NAND2_222(II2415,II2405,II2413);
  nand NAND2_223(WX913,II2414,II2415);
  nand NAND2_224(II2422,WX1001,WX673);
  nand NAND2_225(II2423,WX1001,II2422);
  nand NAND2_226(II2424,WX673,II2422);
  nand NAND2_227(II2421,II2423,II2424);
  nand NAND2_228(II2429,WX737,II2421);
  nand NAND2_229(II2430,WX737,II2429);
  nand NAND2_230(II2431,II2421,II2429);
  nand NAND2_231(II2420,II2430,II2431);
  nand NAND2_232(II2437,WX801,WX865);
  nand NAND2_233(II2438,WX801,II2437);
  nand NAND2_234(II2439,WX865,II2437);
  nand NAND2_235(II2436,II2438,II2439);
  nand NAND2_236(II2444,II2420,II2436);
  nand NAND2_237(II2445,II2420,II2444);
  nand NAND2_238(II2446,II2436,II2444);
  nand NAND2_239(WX914,II2445,II2446);
  nand NAND2_240(II2453,WX1001,WX675);
  nand NAND2_241(II2454,WX1001,II2453);
  nand NAND2_242(II2455,WX675,II2453);
  nand NAND2_243(II2452,II2454,II2455);
  nand NAND2_244(II2460,WX739,II2452);
  nand NAND2_245(II2461,WX739,II2460);
  nand NAND2_246(II2462,II2452,II2460);
  nand NAND2_247(II2451,II2461,II2462);
  nand NAND2_248(II2468,WX803,WX867);
  nand NAND2_249(II2469,WX803,II2468);
  nand NAND2_250(II2470,WX867,II2468);
  nand NAND2_251(II2467,II2469,II2470);
  nand NAND2_252(II2475,II2451,II2467);
  nand NAND2_253(II2476,II2451,II2475);
  nand NAND2_254(II2477,II2467,II2475);
  nand NAND2_255(WX915,II2476,II2477);
  nand NAND2_256(II2484,WX1002,WX677);
  nand NAND2_257(II2485,WX1002,II2484);
  nand NAND2_258(II2486,WX677,II2484);
  nand NAND2_259(II2483,II2485,II2486);
  nand NAND2_260(II2491,WX741,II2483);
  nand NAND2_261(II2492,WX741,II2491);
  nand NAND2_262(II2493,II2483,II2491);
  nand NAND2_263(II2482,II2492,II2493);
  nand NAND2_264(II2499,WX805,WX869);
  nand NAND2_265(II2500,WX805,II2499);
  nand NAND2_266(II2501,WX869,II2499);
  nand NAND2_267(II2498,II2500,II2501);
  nand NAND2_268(II2506,II2482,II2498);
  nand NAND2_269(II2507,II2482,II2506);
  nand NAND2_270(II2508,II2498,II2506);
  nand NAND2_271(WX916,II2507,II2508);
  nand NAND2_272(II2515,WX1002,WX679);
  nand NAND2_273(II2516,WX1002,II2515);
  nand NAND2_274(II2517,WX679,II2515);
  nand NAND2_275(II2514,II2516,II2517);
  nand NAND2_276(II2522,WX743,II2514);
  nand NAND2_277(II2523,WX743,II2522);
  nand NAND2_278(II2524,II2514,II2522);
  nand NAND2_279(II2513,II2523,II2524);
  nand NAND2_280(II2530,WX807,WX871);
  nand NAND2_281(II2531,WX807,II2530);
  nand NAND2_282(II2532,WX871,II2530);
  nand NAND2_283(II2529,II2531,II2532);
  nand NAND2_284(II2537,II2513,II2529);
  nand NAND2_285(II2538,II2513,II2537);
  nand NAND2_286(II2539,II2529,II2537);
  nand NAND2_287(WX917,II2538,II2539);
  nand NAND2_288(II2546,WX1002,WX681);
  nand NAND2_289(II2547,WX1002,II2546);
  nand NAND2_290(II2548,WX681,II2546);
  nand NAND2_291(II2545,II2547,II2548);
  nand NAND2_292(II2553,WX745,II2545);
  nand NAND2_293(II2554,WX745,II2553);
  nand NAND2_294(II2555,II2545,II2553);
  nand NAND2_295(II2544,II2554,II2555);
  nand NAND2_296(II2561,WX809,WX873);
  nand NAND2_297(II2562,WX809,II2561);
  nand NAND2_298(II2563,WX873,II2561);
  nand NAND2_299(II2560,II2562,II2563);
  nand NAND2_300(II2568,II2544,II2560);
  nand NAND2_301(II2569,II2544,II2568);
  nand NAND2_302(II2570,II2560,II2568);
  nand NAND2_303(WX918,II2569,II2570);
  nand NAND2_304(II2577,WX1002,WX683);
  nand NAND2_305(II2578,WX1002,II2577);
  nand NAND2_306(II2579,WX683,II2577);
  nand NAND2_307(II2576,II2578,II2579);
  nand NAND2_308(II2584,WX747,II2576);
  nand NAND2_309(II2585,WX747,II2584);
  nand NAND2_310(II2586,II2576,II2584);
  nand NAND2_311(II2575,II2585,II2586);
  nand NAND2_312(II2592,WX811,WX875);
  nand NAND2_313(II2593,WX811,II2592);
  nand NAND2_314(II2594,WX875,II2592);
  nand NAND2_315(II2591,II2593,II2594);
  nand NAND2_316(II2599,II2575,II2591);
  nand NAND2_317(II2600,II2575,II2599);
  nand NAND2_318(II2601,II2591,II2599);
  nand NAND2_319(WX919,II2600,II2601);
  nand NAND2_320(II2608,WX1002,WX685);
  nand NAND2_321(II2609,WX1002,II2608);
  nand NAND2_322(II2610,WX685,II2608);
  nand NAND2_323(II2607,II2609,II2610);
  nand NAND2_324(II2615,WX749,II2607);
  nand NAND2_325(II2616,WX749,II2615);
  nand NAND2_326(II2617,II2607,II2615);
  nand NAND2_327(II2606,II2616,II2617);
  nand NAND2_328(II2623,WX813,WX877);
  nand NAND2_329(II2624,WX813,II2623);
  nand NAND2_330(II2625,WX877,II2623);
  nand NAND2_331(II2622,II2624,II2625);
  nand NAND2_332(II2630,II2606,II2622);
  nand NAND2_333(II2631,II2606,II2630);
  nand NAND2_334(II2632,II2622,II2630);
  nand NAND2_335(WX920,II2631,II2632);
  nand NAND2_336(II2639,WX1002,WX687);
  nand NAND2_337(II2640,WX1002,II2639);
  nand NAND2_338(II2641,WX687,II2639);
  nand NAND2_339(II2638,II2640,II2641);
  nand NAND2_340(II2646,WX751,II2638);
  nand NAND2_341(II2647,WX751,II2646);
  nand NAND2_342(II2648,II2638,II2646);
  nand NAND2_343(II2637,II2647,II2648);
  nand NAND2_344(II2654,WX815,WX879);
  nand NAND2_345(II2655,WX815,II2654);
  nand NAND2_346(II2656,WX879,II2654);
  nand NAND2_347(II2653,II2655,II2656);
  nand NAND2_348(II2661,II2637,II2653);
  nand NAND2_349(II2662,II2637,II2661);
  nand NAND2_350(II2663,II2653,II2661);
  nand NAND2_351(WX921,II2662,II2663);
  nand NAND2_352(II2670,WX1002,WX689);
  nand NAND2_353(II2671,WX1002,II2670);
  nand NAND2_354(II2672,WX689,II2670);
  nand NAND2_355(II2669,II2671,II2672);
  nand NAND2_356(II2677,WX753,II2669);
  nand NAND2_357(II2678,WX753,II2677);
  nand NAND2_358(II2679,II2669,II2677);
  nand NAND2_359(II2668,II2678,II2679);
  nand NAND2_360(II2685,WX817,WX881);
  nand NAND2_361(II2686,WX817,II2685);
  nand NAND2_362(II2687,WX881,II2685);
  nand NAND2_363(II2684,II2686,II2687);
  nand NAND2_364(II2692,II2668,II2684);
  nand NAND2_365(II2693,II2668,II2692);
  nand NAND2_366(II2694,II2684,II2692);
  nand NAND2_367(WX922,II2693,II2694);
  nand NAND2_368(II2701,WX1002,WX691);
  nand NAND2_369(II2702,WX1002,II2701);
  nand NAND2_370(II2703,WX691,II2701);
  nand NAND2_371(II2700,II2702,II2703);
  nand NAND2_372(II2708,WX755,II2700);
  nand NAND2_373(II2709,WX755,II2708);
  nand NAND2_374(II2710,II2700,II2708);
  nand NAND2_375(II2699,II2709,II2710);
  nand NAND2_376(II2716,WX819,WX883);
  nand NAND2_377(II2717,WX819,II2716);
  nand NAND2_378(II2718,WX883,II2716);
  nand NAND2_379(II2715,II2717,II2718);
  nand NAND2_380(II2723,II2699,II2715);
  nand NAND2_381(II2724,II2699,II2723);
  nand NAND2_382(II2725,II2715,II2723);
  nand NAND2_383(WX923,II2724,II2725);
  nand NAND2_384(II2732,WX1002,WX693);
  nand NAND2_385(II2733,WX1002,II2732);
  nand NAND2_386(II2734,WX693,II2732);
  nand NAND2_387(II2731,II2733,II2734);
  nand NAND2_388(II2739,WX757,II2731);
  nand NAND2_389(II2740,WX757,II2739);
  nand NAND2_390(II2741,II2731,II2739);
  nand NAND2_391(II2730,II2740,II2741);
  nand NAND2_392(II2747,WX821,WX885);
  nand NAND2_393(II2748,WX821,II2747);
  nand NAND2_394(II2749,WX885,II2747);
  nand NAND2_395(II2746,II2748,II2749);
  nand NAND2_396(II2754,II2730,II2746);
  nand NAND2_397(II2755,II2730,II2754);
  nand NAND2_398(II2756,II2746,II2754);
  nand NAND2_399(WX924,II2755,II2756);
  nand NAND2_400(II2763,WX1002,WX695);
  nand NAND2_401(II2764,WX1002,II2763);
  nand NAND2_402(II2765,WX695,II2763);
  nand NAND2_403(II2762,II2764,II2765);
  nand NAND2_404(II2770,WX759,II2762);
  nand NAND2_405(II2771,WX759,II2770);
  nand NAND2_406(II2772,II2762,II2770);
  nand NAND2_407(II2761,II2771,II2772);
  nand NAND2_408(II2778,WX823,WX887);
  nand NAND2_409(II2779,WX823,II2778);
  nand NAND2_410(II2780,WX887,II2778);
  nand NAND2_411(II2777,II2779,II2780);
  nand NAND2_412(II2785,II2761,II2777);
  nand NAND2_413(II2786,II2761,II2785);
  nand NAND2_414(II2787,II2777,II2785);
  nand NAND2_415(WX925,II2786,II2787);
  nand NAND2_416(II2794,WX1002,WX697);
  nand NAND2_417(II2795,WX1002,II2794);
  nand NAND2_418(II2796,WX697,II2794);
  nand NAND2_419(II2793,II2795,II2796);
  nand NAND2_420(II2801,WX761,II2793);
  nand NAND2_421(II2802,WX761,II2801);
  nand NAND2_422(II2803,II2793,II2801);
  nand NAND2_423(II2792,II2802,II2803);
  nand NAND2_424(II2809,WX825,WX889);
  nand NAND2_425(II2810,WX825,II2809);
  nand NAND2_426(II2811,WX889,II2809);
  nand NAND2_427(II2808,II2810,II2811);
  nand NAND2_428(II2816,II2792,II2808);
  nand NAND2_429(II2817,II2792,II2816);
  nand NAND2_430(II2818,II2808,II2816);
  nand NAND2_431(WX926,II2817,II2818);
  nand NAND2_432(II2825,WX1002,WX699);
  nand NAND2_433(II2826,WX1002,II2825);
  nand NAND2_434(II2827,WX699,II2825);
  nand NAND2_435(II2824,II2826,II2827);
  nand NAND2_436(II2832,WX763,II2824);
  nand NAND2_437(II2833,WX763,II2832);
  nand NAND2_438(II2834,II2824,II2832);
  nand NAND2_439(II2823,II2833,II2834);
  nand NAND2_440(II2840,WX827,WX891);
  nand NAND2_441(II2841,WX827,II2840);
  nand NAND2_442(II2842,WX891,II2840);
  nand NAND2_443(II2839,II2841,II2842);
  nand NAND2_444(II2847,II2823,II2839);
  nand NAND2_445(II2848,II2823,II2847);
  nand NAND2_446(II2849,II2839,II2847);
  nand NAND2_447(WX927,II2848,II2849);
  nand NAND2_448(II2856,WX1002,WX701);
  nand NAND2_449(II2857,WX1002,II2856);
  nand NAND2_450(II2858,WX701,II2856);
  nand NAND2_451(II2855,II2857,II2858);
  nand NAND2_452(II2863,WX765,II2855);
  nand NAND2_453(II2864,WX765,II2863);
  nand NAND2_454(II2865,II2855,II2863);
  nand NAND2_455(II2854,II2864,II2865);
  nand NAND2_456(II2871,WX829,WX893);
  nand NAND2_457(II2872,WX829,II2871);
  nand NAND2_458(II2873,WX893,II2871);
  nand NAND2_459(II2870,II2872,II2873);
  nand NAND2_460(II2878,II2854,II2870);
  nand NAND2_461(II2879,II2854,II2878);
  nand NAND2_462(II2880,II2870,II2878);
  nand NAND2_463(WX928,II2879,II2880);
  nand NAND2_464(II2887,WX1002,WX703);
  nand NAND2_465(II2888,WX1002,II2887);
  nand NAND2_466(II2889,WX703,II2887);
  nand NAND2_467(II2886,II2888,II2889);
  nand NAND2_468(II2894,WX767,II2886);
  nand NAND2_469(II2895,WX767,II2894);
  nand NAND2_470(II2896,II2886,II2894);
  nand NAND2_471(II2885,II2895,II2896);
  nand NAND2_472(II2902,WX831,WX895);
  nand NAND2_473(II2903,WX831,II2902);
  nand NAND2_474(II2904,WX895,II2902);
  nand NAND2_475(II2901,II2903,II2904);
  nand NAND2_476(II2909,II2885,II2901);
  nand NAND2_477(II2910,II2885,II2909);
  nand NAND2_478(II2911,II2901,II2909);
  nand NAND2_479(WX929,II2910,II2911);
  nand NAND2_480(II2918,WX1002,WX705);
  nand NAND2_481(II2919,WX1002,II2918);
  nand NAND2_482(II2920,WX705,II2918);
  nand NAND2_483(II2917,II2919,II2920);
  nand NAND2_484(II2925,WX769,II2917);
  nand NAND2_485(II2926,WX769,II2925);
  nand NAND2_486(II2927,II2917,II2925);
  nand NAND2_487(II2916,II2926,II2927);
  nand NAND2_488(II2933,WX833,WX897);
  nand NAND2_489(II2934,WX833,II2933);
  nand NAND2_490(II2935,WX897,II2933);
  nand NAND2_491(II2932,II2934,II2935);
  nand NAND2_492(II2940,II2916,II2932);
  nand NAND2_493(II2941,II2916,II2940);
  nand NAND2_494(II2942,II2932,II2940);
  nand NAND2_495(WX930,II2941,II2942);
  nand NAND2_496(II2949,WX1002,WX707);
  nand NAND2_497(II2950,WX1002,II2949);
  nand NAND2_498(II2951,WX707,II2949);
  nand NAND2_499(II2948,II2950,II2951);
  nand NAND2_500(II2956,WX771,II2948);
  nand NAND2_501(II2957,WX771,II2956);
  nand NAND2_502(II2958,II2948,II2956);
  nand NAND2_503(II2947,II2957,II2958);
  nand NAND2_504(II2964,WX835,WX899);
  nand NAND2_505(II2965,WX835,II2964);
  nand NAND2_506(II2966,WX899,II2964);
  nand NAND2_507(II2963,II2965,II2966);
  nand NAND2_508(II2971,II2947,II2963);
  nand NAND2_509(II2972,II2947,II2971);
  nand NAND2_510(II2973,II2963,II2971);
  nand NAND2_511(WX931,II2972,II2973);
  nand NAND2_512(II3052,WX580,WX485);
  nand NAND2_513(II3053,WX580,II3052);
  nand NAND2_514(II3054,WX485,II3052);
  nand NAND2_515(WX1006,II3053,II3054);
  nand NAND2_516(II3065,WX581,WX487);
  nand NAND2_517(II3066,WX581,II3065);
  nand NAND2_518(II3067,WX487,II3065);
  nand NAND2_519(WX1013,II3066,II3067);
  nand NAND2_520(II3078,WX582,WX489);
  nand NAND2_521(II3079,WX582,II3078);
  nand NAND2_522(II3080,WX489,II3078);
  nand NAND2_523(WX1020,II3079,II3080);
  nand NAND2_524(II3091,WX583,WX491);
  nand NAND2_525(II3092,WX583,II3091);
  nand NAND2_526(II3093,WX491,II3091);
  nand NAND2_527(WX1027,II3092,II3093);
  nand NAND2_528(II3104,WX584,WX493);
  nand NAND2_529(II3105,WX584,II3104);
  nand NAND2_530(II3106,WX493,II3104);
  nand NAND2_531(WX1034,II3105,II3106);
  nand NAND2_532(II3117,WX585,WX495);
  nand NAND2_533(II3118,WX585,II3117);
  nand NAND2_534(II3119,WX495,II3117);
  nand NAND2_535(WX1041,II3118,II3119);
  nand NAND2_536(II3130,WX586,WX497);
  nand NAND2_537(II3131,WX586,II3130);
  nand NAND2_538(II3132,WX497,II3130);
  nand NAND2_539(WX1048,II3131,II3132);
  nand NAND2_540(II3143,WX587,WX499);
  nand NAND2_541(II3144,WX587,II3143);
  nand NAND2_542(II3145,WX499,II3143);
  nand NAND2_543(WX1055,II3144,II3145);
  nand NAND2_544(II3156,WX588,WX501);
  nand NAND2_545(II3157,WX588,II3156);
  nand NAND2_546(II3158,WX501,II3156);
  nand NAND2_547(WX1062,II3157,II3158);
  nand NAND2_548(II3169,WX589,WX503);
  nand NAND2_549(II3170,WX589,II3169);
  nand NAND2_550(II3171,WX503,II3169);
  nand NAND2_551(WX1069,II3170,II3171);
  nand NAND2_552(II3182,WX590,WX505);
  nand NAND2_553(II3183,WX590,II3182);
  nand NAND2_554(II3184,WX505,II3182);
  nand NAND2_555(WX1076,II3183,II3184);
  nand NAND2_556(II3195,WX591,WX507);
  nand NAND2_557(II3196,WX591,II3195);
  nand NAND2_558(II3197,WX507,II3195);
  nand NAND2_559(WX1083,II3196,II3197);
  nand NAND2_560(II3208,WX592,WX509);
  nand NAND2_561(II3209,WX592,II3208);
  nand NAND2_562(II3210,WX509,II3208);
  nand NAND2_563(WX1090,II3209,II3210);
  nand NAND2_564(II3221,WX593,WX511);
  nand NAND2_565(II3222,WX593,II3221);
  nand NAND2_566(II3223,WX511,II3221);
  nand NAND2_567(WX1097,II3222,II3223);
  nand NAND2_568(II3234,WX594,WX513);
  nand NAND2_569(II3235,WX594,II3234);
  nand NAND2_570(II3236,WX513,II3234);
  nand NAND2_571(WX1104,II3235,II3236);
  nand NAND2_572(II3247,WX595,WX515);
  nand NAND2_573(II3248,WX595,II3247);
  nand NAND2_574(II3249,WX515,II3247);
  nand NAND2_575(WX1111,II3248,II3249);
  nand NAND2_576(II3260,WX596,WX517);
  nand NAND2_577(II3261,WX596,II3260);
  nand NAND2_578(II3262,WX517,II3260);
  nand NAND2_579(WX1118,II3261,II3262);
  nand NAND2_580(II3273,WX597,WX519);
  nand NAND2_581(II3274,WX597,II3273);
  nand NAND2_582(II3275,WX519,II3273);
  nand NAND2_583(WX1125,II3274,II3275);
  nand NAND2_584(II3286,WX598,WX521);
  nand NAND2_585(II3287,WX598,II3286);
  nand NAND2_586(II3288,WX521,II3286);
  nand NAND2_587(WX1132,II3287,II3288);
  nand NAND2_588(II3299,WX599,WX523);
  nand NAND2_589(II3300,WX599,II3299);
  nand NAND2_590(II3301,WX523,II3299);
  nand NAND2_591(WX1139,II3300,II3301);
  nand NAND2_592(II3312,WX600,WX525);
  nand NAND2_593(II3313,WX600,II3312);
  nand NAND2_594(II3314,WX525,II3312);
  nand NAND2_595(WX1146,II3313,II3314);
  nand NAND2_596(II3325,WX601,WX527);
  nand NAND2_597(II3326,WX601,II3325);
  nand NAND2_598(II3327,WX527,II3325);
  nand NAND2_599(WX1153,II3326,II3327);
  nand NAND2_600(II3338,WX602,WX529);
  nand NAND2_601(II3339,WX602,II3338);
  nand NAND2_602(II3340,WX529,II3338);
  nand NAND2_603(WX1160,II3339,II3340);
  nand NAND2_604(II3351,WX603,WX531);
  nand NAND2_605(II3352,WX603,II3351);
  nand NAND2_606(II3353,WX531,II3351);
  nand NAND2_607(WX1167,II3352,II3353);
  nand NAND2_608(II3364,WX604,WX533);
  nand NAND2_609(II3365,WX604,II3364);
  nand NAND2_610(II3366,WX533,II3364);
  nand NAND2_611(WX1174,II3365,II3366);
  nand NAND2_612(II3377,WX605,WX535);
  nand NAND2_613(II3378,WX605,II3377);
  nand NAND2_614(II3379,WX535,II3377);
  nand NAND2_615(WX1181,II3378,II3379);
  nand NAND2_616(II3390,WX606,WX537);
  nand NAND2_617(II3391,WX606,II3390);
  nand NAND2_618(II3392,WX537,II3390);
  nand NAND2_619(WX1188,II3391,II3392);
  nand NAND2_620(II3403,WX607,WX539);
  nand NAND2_621(II3404,WX607,II3403);
  nand NAND2_622(II3405,WX539,II3403);
  nand NAND2_623(WX1195,II3404,II3405);
  nand NAND2_624(II3416,WX608,WX541);
  nand NAND2_625(II3417,WX608,II3416);
  nand NAND2_626(II3418,WX541,II3416);
  nand NAND2_627(WX1202,II3417,II3418);
  nand NAND2_628(II3429,WX609,WX543);
  nand NAND2_629(II3430,WX609,II3429);
  nand NAND2_630(II3431,WX543,II3429);
  nand NAND2_631(WX1209,II3430,II3431);
  nand NAND2_632(II3442,WX610,WX545);
  nand NAND2_633(II3443,WX610,II3442);
  nand NAND2_634(II3444,WX545,II3442);
  nand NAND2_635(WX1216,II3443,II3444);
  nand NAND2_636(II3455,WX611,WX547);
  nand NAND2_637(II3456,WX611,II3455);
  nand NAND2_638(II3457,WX547,II3455);
  nand NAND2_639(WX1223,II3456,II3457);
  nand NAND2_640(II3470,WX627,CRC_OUT_9_31);
  nand NAND2_641(II3471,WX627,II3470);
  nand NAND2_642(II3472,CRC_OUT_9_31,II3470);
  nand NAND2_643(II3469,II3471,II3472);
  nand NAND2_644(II3477,CRC_OUT_9_15,II3469);
  nand NAND2_645(II3478,CRC_OUT_9_15,II3477);
  nand NAND2_646(II3479,II3469,II3477);
  nand NAND2_647(WX1231,II3478,II3479);
  nand NAND2_648(II3485,WX632,CRC_OUT_9_31);
  nand NAND2_649(II3486,WX632,II3485);
  nand NAND2_650(II3487,CRC_OUT_9_31,II3485);
  nand NAND2_651(II3484,II3486,II3487);
  nand NAND2_652(II3492,CRC_OUT_9_10,II3484);
  nand NAND2_653(II3493,CRC_OUT_9_10,II3492);
  nand NAND2_654(II3494,II3484,II3492);
  nand NAND2_655(WX1232,II3493,II3494);
  nand NAND2_656(II3500,WX639,CRC_OUT_9_31);
  nand NAND2_657(II3501,WX639,II3500);
  nand NAND2_658(II3502,CRC_OUT_9_31,II3500);
  nand NAND2_659(II3499,II3501,II3502);
  nand NAND2_660(II3507,CRC_OUT_9_3,II3499);
  nand NAND2_661(II3508,CRC_OUT_9_3,II3507);
  nand NAND2_662(II3509,II3499,II3507);
  nand NAND2_663(WX1233,II3508,II3509);
  nand NAND2_664(II3514,WX643,CRC_OUT_9_31);
  nand NAND2_665(II3515,WX643,II3514);
  nand NAND2_666(II3516,CRC_OUT_9_31,II3514);
  nand NAND2_667(WX1234,II3515,II3516);
  nand NAND2_668(II3521,WX612,CRC_OUT_9_30);
  nand NAND2_669(II3522,WX612,II3521);
  nand NAND2_670(II3523,CRC_OUT_9_30,II3521);
  nand NAND2_671(WX1235,II3522,II3523);
  nand NAND2_672(II3528,WX613,CRC_OUT_9_29);
  nand NAND2_673(II3529,WX613,II3528);
  nand NAND2_674(II3530,CRC_OUT_9_29,II3528);
  nand NAND2_675(WX1236,II3529,II3530);
  nand NAND2_676(II3535,WX614,CRC_OUT_9_28);
  nand NAND2_677(II3536,WX614,II3535);
  nand NAND2_678(II3537,CRC_OUT_9_28,II3535);
  nand NAND2_679(WX1237,II3536,II3537);
  nand NAND2_680(II3542,WX615,CRC_OUT_9_27);
  nand NAND2_681(II3543,WX615,II3542);
  nand NAND2_682(II3544,CRC_OUT_9_27,II3542);
  nand NAND2_683(WX1238,II3543,II3544);
  nand NAND2_684(II3549,WX616,CRC_OUT_9_26);
  nand NAND2_685(II3550,WX616,II3549);
  nand NAND2_686(II3551,CRC_OUT_9_26,II3549);
  nand NAND2_687(WX1239,II3550,II3551);
  nand NAND2_688(II3556,WX617,CRC_OUT_9_25);
  nand NAND2_689(II3557,WX617,II3556);
  nand NAND2_690(II3558,CRC_OUT_9_25,II3556);
  nand NAND2_691(WX1240,II3557,II3558);
  nand NAND2_692(II3563,WX618,CRC_OUT_9_24);
  nand NAND2_693(II3564,WX618,II3563);
  nand NAND2_694(II3565,CRC_OUT_9_24,II3563);
  nand NAND2_695(WX1241,II3564,II3565);
  nand NAND2_696(II3570,WX619,CRC_OUT_9_23);
  nand NAND2_697(II3571,WX619,II3570);
  nand NAND2_698(II3572,CRC_OUT_9_23,II3570);
  nand NAND2_699(WX1242,II3571,II3572);
  nand NAND2_700(II3577,WX620,CRC_OUT_9_22);
  nand NAND2_701(II3578,WX620,II3577);
  nand NAND2_702(II3579,CRC_OUT_9_22,II3577);
  nand NAND2_703(WX1243,II3578,II3579);
  nand NAND2_704(II3584,WX621,CRC_OUT_9_21);
  nand NAND2_705(II3585,WX621,II3584);
  nand NAND2_706(II3586,CRC_OUT_9_21,II3584);
  nand NAND2_707(WX1244,II3585,II3586);
  nand NAND2_708(II3591,WX622,CRC_OUT_9_20);
  nand NAND2_709(II3592,WX622,II3591);
  nand NAND2_710(II3593,CRC_OUT_9_20,II3591);
  nand NAND2_711(WX1245,II3592,II3593);
  nand NAND2_712(II3598,WX623,CRC_OUT_9_19);
  nand NAND2_713(II3599,WX623,II3598);
  nand NAND2_714(II3600,CRC_OUT_9_19,II3598);
  nand NAND2_715(WX1246,II3599,II3600);
  nand NAND2_716(II3605,WX624,CRC_OUT_9_18);
  nand NAND2_717(II3606,WX624,II3605);
  nand NAND2_718(II3607,CRC_OUT_9_18,II3605);
  nand NAND2_719(WX1247,II3606,II3607);
  nand NAND2_720(II3612,WX625,CRC_OUT_9_17);
  nand NAND2_721(II3613,WX625,II3612);
  nand NAND2_722(II3614,CRC_OUT_9_17,II3612);
  nand NAND2_723(WX1248,II3613,II3614);
  nand NAND2_724(II3619,WX626,CRC_OUT_9_16);
  nand NAND2_725(II3620,WX626,II3619);
  nand NAND2_726(II3621,CRC_OUT_9_16,II3619);
  nand NAND2_727(WX1249,II3620,II3621);
  nand NAND2_728(II3626,WX628,CRC_OUT_9_14);
  nand NAND2_729(II3627,WX628,II3626);
  nand NAND2_730(II3628,CRC_OUT_9_14,II3626);
  nand NAND2_731(WX1250,II3627,II3628);
  nand NAND2_732(II3633,WX629,CRC_OUT_9_13);
  nand NAND2_733(II3634,WX629,II3633);
  nand NAND2_734(II3635,CRC_OUT_9_13,II3633);
  nand NAND2_735(WX1251,II3634,II3635);
  nand NAND2_736(II3640,WX630,CRC_OUT_9_12);
  nand NAND2_737(II3641,WX630,II3640);
  nand NAND2_738(II3642,CRC_OUT_9_12,II3640);
  nand NAND2_739(WX1252,II3641,II3642);
  nand NAND2_740(II3647,WX631,CRC_OUT_9_11);
  nand NAND2_741(II3648,WX631,II3647);
  nand NAND2_742(II3649,CRC_OUT_9_11,II3647);
  nand NAND2_743(WX1253,II3648,II3649);
  nand NAND2_744(II3654,WX633,CRC_OUT_9_9);
  nand NAND2_745(II3655,WX633,II3654);
  nand NAND2_746(II3656,CRC_OUT_9_9,II3654);
  nand NAND2_747(WX1254,II3655,II3656);
  nand NAND2_748(II3661,WX634,CRC_OUT_9_8);
  nand NAND2_749(II3662,WX634,II3661);
  nand NAND2_750(II3663,CRC_OUT_9_8,II3661);
  nand NAND2_751(WX1255,II3662,II3663);
  nand NAND2_752(II3668,WX635,CRC_OUT_9_7);
  nand NAND2_753(II3669,WX635,II3668);
  nand NAND2_754(II3670,CRC_OUT_9_7,II3668);
  nand NAND2_755(WX1256,II3669,II3670);
  nand NAND2_756(II3675,WX636,CRC_OUT_9_6);
  nand NAND2_757(II3676,WX636,II3675);
  nand NAND2_758(II3677,CRC_OUT_9_6,II3675);
  nand NAND2_759(WX1257,II3676,II3677);
  nand NAND2_760(II3682,WX637,CRC_OUT_9_5);
  nand NAND2_761(II3683,WX637,II3682);
  nand NAND2_762(II3684,CRC_OUT_9_5,II3682);
  nand NAND2_763(WX1258,II3683,II3684);
  nand NAND2_764(II3689,WX638,CRC_OUT_9_4);
  nand NAND2_765(II3690,WX638,II3689);
  nand NAND2_766(II3691,CRC_OUT_9_4,II3689);
  nand NAND2_767(WX1259,II3690,II3691);
  nand NAND2_768(II3696,WX640,CRC_OUT_9_2);
  nand NAND2_769(II3697,WX640,II3696);
  nand NAND2_770(II3698,CRC_OUT_9_2,II3696);
  nand NAND2_771(WX1260,II3697,II3698);
  nand NAND2_772(II3703,WX641,CRC_OUT_9_1);
  nand NAND2_773(II3704,WX641,II3703);
  nand NAND2_774(II3705,CRC_OUT_9_1,II3703);
  nand NAND2_775(WX1261,II3704,II3705);
  nand NAND2_776(II3710,WX642,CRC_OUT_9_0);
  nand NAND2_777(II3711,WX642,II3710);
  nand NAND2_778(II3712,CRC_OUT_9_0,II3710);
  nand NAND2_779(WX1262,II3711,II3712);
  nand NAND2_780(II5993,WX2294,WX1938);
  nand NAND2_781(II5994,WX2294,II5993);
  nand NAND2_782(II5995,WX1938,II5993);
  nand NAND2_783(II5992,II5994,II5995);
  nand NAND2_784(II6000,WX2002,II5992);
  nand NAND2_785(II6001,WX2002,II6000);
  nand NAND2_786(II6002,II5992,II6000);
  nand NAND2_787(II5991,II6001,II6002);
  nand NAND2_788(II6008,WX2066,WX2130);
  nand NAND2_789(II6009,WX2066,II6008);
  nand NAND2_790(II6010,WX2130,II6008);
  nand NAND2_791(II6007,II6009,II6010);
  nand NAND2_792(II6015,II5991,II6007);
  nand NAND2_793(II6016,II5991,II6015);
  nand NAND2_794(II6017,II6007,II6015);
  nand NAND2_795(WX2193,II6016,II6017);
  nand NAND2_796(II6024,WX2294,WX1940);
  nand NAND2_797(II6025,WX2294,II6024);
  nand NAND2_798(II6026,WX1940,II6024);
  nand NAND2_799(II6023,II6025,II6026);
  nand NAND2_800(II6031,WX2004,II6023);
  nand NAND2_801(II6032,WX2004,II6031);
  nand NAND2_802(II6033,II6023,II6031);
  nand NAND2_803(II6022,II6032,II6033);
  nand NAND2_804(II6039,WX2068,WX2132);
  nand NAND2_805(II6040,WX2068,II6039);
  nand NAND2_806(II6041,WX2132,II6039);
  nand NAND2_807(II6038,II6040,II6041);
  nand NAND2_808(II6046,II6022,II6038);
  nand NAND2_809(II6047,II6022,II6046);
  nand NAND2_810(II6048,II6038,II6046);
  nand NAND2_811(WX2194,II6047,II6048);
  nand NAND2_812(II6055,WX2294,WX1942);
  nand NAND2_813(II6056,WX2294,II6055);
  nand NAND2_814(II6057,WX1942,II6055);
  nand NAND2_815(II6054,II6056,II6057);
  nand NAND2_816(II6062,WX2006,II6054);
  nand NAND2_817(II6063,WX2006,II6062);
  nand NAND2_818(II6064,II6054,II6062);
  nand NAND2_819(II6053,II6063,II6064);
  nand NAND2_820(II6070,WX2070,WX2134);
  nand NAND2_821(II6071,WX2070,II6070);
  nand NAND2_822(II6072,WX2134,II6070);
  nand NAND2_823(II6069,II6071,II6072);
  nand NAND2_824(II6077,II6053,II6069);
  nand NAND2_825(II6078,II6053,II6077);
  nand NAND2_826(II6079,II6069,II6077);
  nand NAND2_827(WX2195,II6078,II6079);
  nand NAND2_828(II6086,WX2294,WX1944);
  nand NAND2_829(II6087,WX2294,II6086);
  nand NAND2_830(II6088,WX1944,II6086);
  nand NAND2_831(II6085,II6087,II6088);
  nand NAND2_832(II6093,WX2008,II6085);
  nand NAND2_833(II6094,WX2008,II6093);
  nand NAND2_834(II6095,II6085,II6093);
  nand NAND2_835(II6084,II6094,II6095);
  nand NAND2_836(II6101,WX2072,WX2136);
  nand NAND2_837(II6102,WX2072,II6101);
  nand NAND2_838(II6103,WX2136,II6101);
  nand NAND2_839(II6100,II6102,II6103);
  nand NAND2_840(II6108,II6084,II6100);
  nand NAND2_841(II6109,II6084,II6108);
  nand NAND2_842(II6110,II6100,II6108);
  nand NAND2_843(WX2196,II6109,II6110);
  nand NAND2_844(II6117,WX2294,WX1946);
  nand NAND2_845(II6118,WX2294,II6117);
  nand NAND2_846(II6119,WX1946,II6117);
  nand NAND2_847(II6116,II6118,II6119);
  nand NAND2_848(II6124,WX2010,II6116);
  nand NAND2_849(II6125,WX2010,II6124);
  nand NAND2_850(II6126,II6116,II6124);
  nand NAND2_851(II6115,II6125,II6126);
  nand NAND2_852(II6132,WX2074,WX2138);
  nand NAND2_853(II6133,WX2074,II6132);
  nand NAND2_854(II6134,WX2138,II6132);
  nand NAND2_855(II6131,II6133,II6134);
  nand NAND2_856(II6139,II6115,II6131);
  nand NAND2_857(II6140,II6115,II6139);
  nand NAND2_858(II6141,II6131,II6139);
  nand NAND2_859(WX2197,II6140,II6141);
  nand NAND2_860(II6148,WX2294,WX1948);
  nand NAND2_861(II6149,WX2294,II6148);
  nand NAND2_862(II6150,WX1948,II6148);
  nand NAND2_863(II6147,II6149,II6150);
  nand NAND2_864(II6155,WX2012,II6147);
  nand NAND2_865(II6156,WX2012,II6155);
  nand NAND2_866(II6157,II6147,II6155);
  nand NAND2_867(II6146,II6156,II6157);
  nand NAND2_868(II6163,WX2076,WX2140);
  nand NAND2_869(II6164,WX2076,II6163);
  nand NAND2_870(II6165,WX2140,II6163);
  nand NAND2_871(II6162,II6164,II6165);
  nand NAND2_872(II6170,II6146,II6162);
  nand NAND2_873(II6171,II6146,II6170);
  nand NAND2_874(II6172,II6162,II6170);
  nand NAND2_875(WX2198,II6171,II6172);
  nand NAND2_876(II6179,WX2294,WX1950);
  nand NAND2_877(II6180,WX2294,II6179);
  nand NAND2_878(II6181,WX1950,II6179);
  nand NAND2_879(II6178,II6180,II6181);
  nand NAND2_880(II6186,WX2014,II6178);
  nand NAND2_881(II6187,WX2014,II6186);
  nand NAND2_882(II6188,II6178,II6186);
  nand NAND2_883(II6177,II6187,II6188);
  nand NAND2_884(II6194,WX2078,WX2142);
  nand NAND2_885(II6195,WX2078,II6194);
  nand NAND2_886(II6196,WX2142,II6194);
  nand NAND2_887(II6193,II6195,II6196);
  nand NAND2_888(II6201,II6177,II6193);
  nand NAND2_889(II6202,II6177,II6201);
  nand NAND2_890(II6203,II6193,II6201);
  nand NAND2_891(WX2199,II6202,II6203);
  nand NAND2_892(II6210,WX2294,WX1952);
  nand NAND2_893(II6211,WX2294,II6210);
  nand NAND2_894(II6212,WX1952,II6210);
  nand NAND2_895(II6209,II6211,II6212);
  nand NAND2_896(II6217,WX2016,II6209);
  nand NAND2_897(II6218,WX2016,II6217);
  nand NAND2_898(II6219,II6209,II6217);
  nand NAND2_899(II6208,II6218,II6219);
  nand NAND2_900(II6225,WX2080,WX2144);
  nand NAND2_901(II6226,WX2080,II6225);
  nand NAND2_902(II6227,WX2144,II6225);
  nand NAND2_903(II6224,II6226,II6227);
  nand NAND2_904(II6232,II6208,II6224);
  nand NAND2_905(II6233,II6208,II6232);
  nand NAND2_906(II6234,II6224,II6232);
  nand NAND2_907(WX2200,II6233,II6234);
  nand NAND2_908(II6241,WX2294,WX1954);
  nand NAND2_909(II6242,WX2294,II6241);
  nand NAND2_910(II6243,WX1954,II6241);
  nand NAND2_911(II6240,II6242,II6243);
  nand NAND2_912(II6248,WX2018,II6240);
  nand NAND2_913(II6249,WX2018,II6248);
  nand NAND2_914(II6250,II6240,II6248);
  nand NAND2_915(II6239,II6249,II6250);
  nand NAND2_916(II6256,WX2082,WX2146);
  nand NAND2_917(II6257,WX2082,II6256);
  nand NAND2_918(II6258,WX2146,II6256);
  nand NAND2_919(II6255,II6257,II6258);
  nand NAND2_920(II6263,II6239,II6255);
  nand NAND2_921(II6264,II6239,II6263);
  nand NAND2_922(II6265,II6255,II6263);
  nand NAND2_923(WX2201,II6264,II6265);
  nand NAND2_924(II6272,WX2294,WX1956);
  nand NAND2_925(II6273,WX2294,II6272);
  nand NAND2_926(II6274,WX1956,II6272);
  nand NAND2_927(II6271,II6273,II6274);
  nand NAND2_928(II6279,WX2020,II6271);
  nand NAND2_929(II6280,WX2020,II6279);
  nand NAND2_930(II6281,II6271,II6279);
  nand NAND2_931(II6270,II6280,II6281);
  nand NAND2_932(II6287,WX2084,WX2148);
  nand NAND2_933(II6288,WX2084,II6287);
  nand NAND2_934(II6289,WX2148,II6287);
  nand NAND2_935(II6286,II6288,II6289);
  nand NAND2_936(II6294,II6270,II6286);
  nand NAND2_937(II6295,II6270,II6294);
  nand NAND2_938(II6296,II6286,II6294);
  nand NAND2_939(WX2202,II6295,II6296);
  nand NAND2_940(II6303,WX2294,WX1958);
  nand NAND2_941(II6304,WX2294,II6303);
  nand NAND2_942(II6305,WX1958,II6303);
  nand NAND2_943(II6302,II6304,II6305);
  nand NAND2_944(II6310,WX2022,II6302);
  nand NAND2_945(II6311,WX2022,II6310);
  nand NAND2_946(II6312,II6302,II6310);
  nand NAND2_947(II6301,II6311,II6312);
  nand NAND2_948(II6318,WX2086,WX2150);
  nand NAND2_949(II6319,WX2086,II6318);
  nand NAND2_950(II6320,WX2150,II6318);
  nand NAND2_951(II6317,II6319,II6320);
  nand NAND2_952(II6325,II6301,II6317);
  nand NAND2_953(II6326,II6301,II6325);
  nand NAND2_954(II6327,II6317,II6325);
  nand NAND2_955(WX2203,II6326,II6327);
  nand NAND2_956(II6334,WX2294,WX1960);
  nand NAND2_957(II6335,WX2294,II6334);
  nand NAND2_958(II6336,WX1960,II6334);
  nand NAND2_959(II6333,II6335,II6336);
  nand NAND2_960(II6341,WX2024,II6333);
  nand NAND2_961(II6342,WX2024,II6341);
  nand NAND2_962(II6343,II6333,II6341);
  nand NAND2_963(II6332,II6342,II6343);
  nand NAND2_964(II6349,WX2088,WX2152);
  nand NAND2_965(II6350,WX2088,II6349);
  nand NAND2_966(II6351,WX2152,II6349);
  nand NAND2_967(II6348,II6350,II6351);
  nand NAND2_968(II6356,II6332,II6348);
  nand NAND2_969(II6357,II6332,II6356);
  nand NAND2_970(II6358,II6348,II6356);
  nand NAND2_971(WX2204,II6357,II6358);
  nand NAND2_972(II6365,WX2294,WX1962);
  nand NAND2_973(II6366,WX2294,II6365);
  nand NAND2_974(II6367,WX1962,II6365);
  nand NAND2_975(II6364,II6366,II6367);
  nand NAND2_976(II6372,WX2026,II6364);
  nand NAND2_977(II6373,WX2026,II6372);
  nand NAND2_978(II6374,II6364,II6372);
  nand NAND2_979(II6363,II6373,II6374);
  nand NAND2_980(II6380,WX2090,WX2154);
  nand NAND2_981(II6381,WX2090,II6380);
  nand NAND2_982(II6382,WX2154,II6380);
  nand NAND2_983(II6379,II6381,II6382);
  nand NAND2_984(II6387,II6363,II6379);
  nand NAND2_985(II6388,II6363,II6387);
  nand NAND2_986(II6389,II6379,II6387);
  nand NAND2_987(WX2205,II6388,II6389);
  nand NAND2_988(II6396,WX2294,WX1964);
  nand NAND2_989(II6397,WX2294,II6396);
  nand NAND2_990(II6398,WX1964,II6396);
  nand NAND2_991(II6395,II6397,II6398);
  nand NAND2_992(II6403,WX2028,II6395);
  nand NAND2_993(II6404,WX2028,II6403);
  nand NAND2_994(II6405,II6395,II6403);
  nand NAND2_995(II6394,II6404,II6405);
  nand NAND2_996(II6411,WX2092,WX2156);
  nand NAND2_997(II6412,WX2092,II6411);
  nand NAND2_998(II6413,WX2156,II6411);
  nand NAND2_999(II6410,II6412,II6413);
  nand NAND2_1000(II6418,II6394,II6410);
  nand NAND2_1001(II6419,II6394,II6418);
  nand NAND2_1002(II6420,II6410,II6418);
  nand NAND2_1003(WX2206,II6419,II6420);
  nand NAND2_1004(II6427,WX2294,WX1966);
  nand NAND2_1005(II6428,WX2294,II6427);
  nand NAND2_1006(II6429,WX1966,II6427);
  nand NAND2_1007(II6426,II6428,II6429);
  nand NAND2_1008(II6434,WX2030,II6426);
  nand NAND2_1009(II6435,WX2030,II6434);
  nand NAND2_1010(II6436,II6426,II6434);
  nand NAND2_1011(II6425,II6435,II6436);
  nand NAND2_1012(II6442,WX2094,WX2158);
  nand NAND2_1013(II6443,WX2094,II6442);
  nand NAND2_1014(II6444,WX2158,II6442);
  nand NAND2_1015(II6441,II6443,II6444);
  nand NAND2_1016(II6449,II6425,II6441);
  nand NAND2_1017(II6450,II6425,II6449);
  nand NAND2_1018(II6451,II6441,II6449);
  nand NAND2_1019(WX2207,II6450,II6451);
  nand NAND2_1020(II6458,WX2294,WX1968);
  nand NAND2_1021(II6459,WX2294,II6458);
  nand NAND2_1022(II6460,WX1968,II6458);
  nand NAND2_1023(II6457,II6459,II6460);
  nand NAND2_1024(II6465,WX2032,II6457);
  nand NAND2_1025(II6466,WX2032,II6465);
  nand NAND2_1026(II6467,II6457,II6465);
  nand NAND2_1027(II6456,II6466,II6467);
  nand NAND2_1028(II6473,WX2096,WX2160);
  nand NAND2_1029(II6474,WX2096,II6473);
  nand NAND2_1030(II6475,WX2160,II6473);
  nand NAND2_1031(II6472,II6474,II6475);
  nand NAND2_1032(II6480,II6456,II6472);
  nand NAND2_1033(II6481,II6456,II6480);
  nand NAND2_1034(II6482,II6472,II6480);
  nand NAND2_1035(WX2208,II6481,II6482);
  nand NAND2_1036(II6489,WX2295,WX1970);
  nand NAND2_1037(II6490,WX2295,II6489);
  nand NAND2_1038(II6491,WX1970,II6489);
  nand NAND2_1039(II6488,II6490,II6491);
  nand NAND2_1040(II6496,WX2034,II6488);
  nand NAND2_1041(II6497,WX2034,II6496);
  nand NAND2_1042(II6498,II6488,II6496);
  nand NAND2_1043(II6487,II6497,II6498);
  nand NAND2_1044(II6504,WX2098,WX2162);
  nand NAND2_1045(II6505,WX2098,II6504);
  nand NAND2_1046(II6506,WX2162,II6504);
  nand NAND2_1047(II6503,II6505,II6506);
  nand NAND2_1048(II6511,II6487,II6503);
  nand NAND2_1049(II6512,II6487,II6511);
  nand NAND2_1050(II6513,II6503,II6511);
  nand NAND2_1051(WX2209,II6512,II6513);
  nand NAND2_1052(II6520,WX2295,WX1972);
  nand NAND2_1053(II6521,WX2295,II6520);
  nand NAND2_1054(II6522,WX1972,II6520);
  nand NAND2_1055(II6519,II6521,II6522);
  nand NAND2_1056(II6527,WX2036,II6519);
  nand NAND2_1057(II6528,WX2036,II6527);
  nand NAND2_1058(II6529,II6519,II6527);
  nand NAND2_1059(II6518,II6528,II6529);
  nand NAND2_1060(II6535,WX2100,WX2164);
  nand NAND2_1061(II6536,WX2100,II6535);
  nand NAND2_1062(II6537,WX2164,II6535);
  nand NAND2_1063(II6534,II6536,II6537);
  nand NAND2_1064(II6542,II6518,II6534);
  nand NAND2_1065(II6543,II6518,II6542);
  nand NAND2_1066(II6544,II6534,II6542);
  nand NAND2_1067(WX2210,II6543,II6544);
  nand NAND2_1068(II6551,WX2295,WX1974);
  nand NAND2_1069(II6552,WX2295,II6551);
  nand NAND2_1070(II6553,WX1974,II6551);
  nand NAND2_1071(II6550,II6552,II6553);
  nand NAND2_1072(II6558,WX2038,II6550);
  nand NAND2_1073(II6559,WX2038,II6558);
  nand NAND2_1074(II6560,II6550,II6558);
  nand NAND2_1075(II6549,II6559,II6560);
  nand NAND2_1076(II6566,WX2102,WX2166);
  nand NAND2_1077(II6567,WX2102,II6566);
  nand NAND2_1078(II6568,WX2166,II6566);
  nand NAND2_1079(II6565,II6567,II6568);
  nand NAND2_1080(II6573,II6549,II6565);
  nand NAND2_1081(II6574,II6549,II6573);
  nand NAND2_1082(II6575,II6565,II6573);
  nand NAND2_1083(WX2211,II6574,II6575);
  nand NAND2_1084(II6582,WX2295,WX1976);
  nand NAND2_1085(II6583,WX2295,II6582);
  nand NAND2_1086(II6584,WX1976,II6582);
  nand NAND2_1087(II6581,II6583,II6584);
  nand NAND2_1088(II6589,WX2040,II6581);
  nand NAND2_1089(II6590,WX2040,II6589);
  nand NAND2_1090(II6591,II6581,II6589);
  nand NAND2_1091(II6580,II6590,II6591);
  nand NAND2_1092(II6597,WX2104,WX2168);
  nand NAND2_1093(II6598,WX2104,II6597);
  nand NAND2_1094(II6599,WX2168,II6597);
  nand NAND2_1095(II6596,II6598,II6599);
  nand NAND2_1096(II6604,II6580,II6596);
  nand NAND2_1097(II6605,II6580,II6604);
  nand NAND2_1098(II6606,II6596,II6604);
  nand NAND2_1099(WX2212,II6605,II6606);
  nand NAND2_1100(II6613,WX2295,WX1978);
  nand NAND2_1101(II6614,WX2295,II6613);
  nand NAND2_1102(II6615,WX1978,II6613);
  nand NAND2_1103(II6612,II6614,II6615);
  nand NAND2_1104(II6620,WX2042,II6612);
  nand NAND2_1105(II6621,WX2042,II6620);
  nand NAND2_1106(II6622,II6612,II6620);
  nand NAND2_1107(II6611,II6621,II6622);
  nand NAND2_1108(II6628,WX2106,WX2170);
  nand NAND2_1109(II6629,WX2106,II6628);
  nand NAND2_1110(II6630,WX2170,II6628);
  nand NAND2_1111(II6627,II6629,II6630);
  nand NAND2_1112(II6635,II6611,II6627);
  nand NAND2_1113(II6636,II6611,II6635);
  nand NAND2_1114(II6637,II6627,II6635);
  nand NAND2_1115(WX2213,II6636,II6637);
  nand NAND2_1116(II6644,WX2295,WX1980);
  nand NAND2_1117(II6645,WX2295,II6644);
  nand NAND2_1118(II6646,WX1980,II6644);
  nand NAND2_1119(II6643,II6645,II6646);
  nand NAND2_1120(II6651,WX2044,II6643);
  nand NAND2_1121(II6652,WX2044,II6651);
  nand NAND2_1122(II6653,II6643,II6651);
  nand NAND2_1123(II6642,II6652,II6653);
  nand NAND2_1124(II6659,WX2108,WX2172);
  nand NAND2_1125(II6660,WX2108,II6659);
  nand NAND2_1126(II6661,WX2172,II6659);
  nand NAND2_1127(II6658,II6660,II6661);
  nand NAND2_1128(II6666,II6642,II6658);
  nand NAND2_1129(II6667,II6642,II6666);
  nand NAND2_1130(II6668,II6658,II6666);
  nand NAND2_1131(WX2214,II6667,II6668);
  nand NAND2_1132(II6675,WX2295,WX1982);
  nand NAND2_1133(II6676,WX2295,II6675);
  nand NAND2_1134(II6677,WX1982,II6675);
  nand NAND2_1135(II6674,II6676,II6677);
  nand NAND2_1136(II6682,WX2046,II6674);
  nand NAND2_1137(II6683,WX2046,II6682);
  nand NAND2_1138(II6684,II6674,II6682);
  nand NAND2_1139(II6673,II6683,II6684);
  nand NAND2_1140(II6690,WX2110,WX2174);
  nand NAND2_1141(II6691,WX2110,II6690);
  nand NAND2_1142(II6692,WX2174,II6690);
  nand NAND2_1143(II6689,II6691,II6692);
  nand NAND2_1144(II6697,II6673,II6689);
  nand NAND2_1145(II6698,II6673,II6697);
  nand NAND2_1146(II6699,II6689,II6697);
  nand NAND2_1147(WX2215,II6698,II6699);
  nand NAND2_1148(II6706,WX2295,WX1984);
  nand NAND2_1149(II6707,WX2295,II6706);
  nand NAND2_1150(II6708,WX1984,II6706);
  nand NAND2_1151(II6705,II6707,II6708);
  nand NAND2_1152(II6713,WX2048,II6705);
  nand NAND2_1153(II6714,WX2048,II6713);
  nand NAND2_1154(II6715,II6705,II6713);
  nand NAND2_1155(II6704,II6714,II6715);
  nand NAND2_1156(II6721,WX2112,WX2176);
  nand NAND2_1157(II6722,WX2112,II6721);
  nand NAND2_1158(II6723,WX2176,II6721);
  nand NAND2_1159(II6720,II6722,II6723);
  nand NAND2_1160(II6728,II6704,II6720);
  nand NAND2_1161(II6729,II6704,II6728);
  nand NAND2_1162(II6730,II6720,II6728);
  nand NAND2_1163(WX2216,II6729,II6730);
  nand NAND2_1164(II6737,WX2295,WX1986);
  nand NAND2_1165(II6738,WX2295,II6737);
  nand NAND2_1166(II6739,WX1986,II6737);
  nand NAND2_1167(II6736,II6738,II6739);
  nand NAND2_1168(II6744,WX2050,II6736);
  nand NAND2_1169(II6745,WX2050,II6744);
  nand NAND2_1170(II6746,II6736,II6744);
  nand NAND2_1171(II6735,II6745,II6746);
  nand NAND2_1172(II6752,WX2114,WX2178);
  nand NAND2_1173(II6753,WX2114,II6752);
  nand NAND2_1174(II6754,WX2178,II6752);
  nand NAND2_1175(II6751,II6753,II6754);
  nand NAND2_1176(II6759,II6735,II6751);
  nand NAND2_1177(II6760,II6735,II6759);
  nand NAND2_1178(II6761,II6751,II6759);
  nand NAND2_1179(WX2217,II6760,II6761);
  nand NAND2_1180(II6768,WX2295,WX1988);
  nand NAND2_1181(II6769,WX2295,II6768);
  nand NAND2_1182(II6770,WX1988,II6768);
  nand NAND2_1183(II6767,II6769,II6770);
  nand NAND2_1184(II6775,WX2052,II6767);
  nand NAND2_1185(II6776,WX2052,II6775);
  nand NAND2_1186(II6777,II6767,II6775);
  nand NAND2_1187(II6766,II6776,II6777);
  nand NAND2_1188(II6783,WX2116,WX2180);
  nand NAND2_1189(II6784,WX2116,II6783);
  nand NAND2_1190(II6785,WX2180,II6783);
  nand NAND2_1191(II6782,II6784,II6785);
  nand NAND2_1192(II6790,II6766,II6782);
  nand NAND2_1193(II6791,II6766,II6790);
  nand NAND2_1194(II6792,II6782,II6790);
  nand NAND2_1195(WX2218,II6791,II6792);
  nand NAND2_1196(II6799,WX2295,WX1990);
  nand NAND2_1197(II6800,WX2295,II6799);
  nand NAND2_1198(II6801,WX1990,II6799);
  nand NAND2_1199(II6798,II6800,II6801);
  nand NAND2_1200(II6806,WX2054,II6798);
  nand NAND2_1201(II6807,WX2054,II6806);
  nand NAND2_1202(II6808,II6798,II6806);
  nand NAND2_1203(II6797,II6807,II6808);
  nand NAND2_1204(II6814,WX2118,WX2182);
  nand NAND2_1205(II6815,WX2118,II6814);
  nand NAND2_1206(II6816,WX2182,II6814);
  nand NAND2_1207(II6813,II6815,II6816);
  nand NAND2_1208(II6821,II6797,II6813);
  nand NAND2_1209(II6822,II6797,II6821);
  nand NAND2_1210(II6823,II6813,II6821);
  nand NAND2_1211(WX2219,II6822,II6823);
  nand NAND2_1212(II6830,WX2295,WX1992);
  nand NAND2_1213(II6831,WX2295,II6830);
  nand NAND2_1214(II6832,WX1992,II6830);
  nand NAND2_1215(II6829,II6831,II6832);
  nand NAND2_1216(II6837,WX2056,II6829);
  nand NAND2_1217(II6838,WX2056,II6837);
  nand NAND2_1218(II6839,II6829,II6837);
  nand NAND2_1219(II6828,II6838,II6839);
  nand NAND2_1220(II6845,WX2120,WX2184);
  nand NAND2_1221(II6846,WX2120,II6845);
  nand NAND2_1222(II6847,WX2184,II6845);
  nand NAND2_1223(II6844,II6846,II6847);
  nand NAND2_1224(II6852,II6828,II6844);
  nand NAND2_1225(II6853,II6828,II6852);
  nand NAND2_1226(II6854,II6844,II6852);
  nand NAND2_1227(WX2220,II6853,II6854);
  nand NAND2_1228(II6861,WX2295,WX1994);
  nand NAND2_1229(II6862,WX2295,II6861);
  nand NAND2_1230(II6863,WX1994,II6861);
  nand NAND2_1231(II6860,II6862,II6863);
  nand NAND2_1232(II6868,WX2058,II6860);
  nand NAND2_1233(II6869,WX2058,II6868);
  nand NAND2_1234(II6870,II6860,II6868);
  nand NAND2_1235(II6859,II6869,II6870);
  nand NAND2_1236(II6876,WX2122,WX2186);
  nand NAND2_1237(II6877,WX2122,II6876);
  nand NAND2_1238(II6878,WX2186,II6876);
  nand NAND2_1239(II6875,II6877,II6878);
  nand NAND2_1240(II6883,II6859,II6875);
  nand NAND2_1241(II6884,II6859,II6883);
  nand NAND2_1242(II6885,II6875,II6883);
  nand NAND2_1243(WX2221,II6884,II6885);
  nand NAND2_1244(II6892,WX2295,WX1996);
  nand NAND2_1245(II6893,WX2295,II6892);
  nand NAND2_1246(II6894,WX1996,II6892);
  nand NAND2_1247(II6891,II6893,II6894);
  nand NAND2_1248(II6899,WX2060,II6891);
  nand NAND2_1249(II6900,WX2060,II6899);
  nand NAND2_1250(II6901,II6891,II6899);
  nand NAND2_1251(II6890,II6900,II6901);
  nand NAND2_1252(II6907,WX2124,WX2188);
  nand NAND2_1253(II6908,WX2124,II6907);
  nand NAND2_1254(II6909,WX2188,II6907);
  nand NAND2_1255(II6906,II6908,II6909);
  nand NAND2_1256(II6914,II6890,II6906);
  nand NAND2_1257(II6915,II6890,II6914);
  nand NAND2_1258(II6916,II6906,II6914);
  nand NAND2_1259(WX2222,II6915,II6916);
  nand NAND2_1260(II6923,WX2295,WX1998);
  nand NAND2_1261(II6924,WX2295,II6923);
  nand NAND2_1262(II6925,WX1998,II6923);
  nand NAND2_1263(II6922,II6924,II6925);
  nand NAND2_1264(II6930,WX2062,II6922);
  nand NAND2_1265(II6931,WX2062,II6930);
  nand NAND2_1266(II6932,II6922,II6930);
  nand NAND2_1267(II6921,II6931,II6932);
  nand NAND2_1268(II6938,WX2126,WX2190);
  nand NAND2_1269(II6939,WX2126,II6938);
  nand NAND2_1270(II6940,WX2190,II6938);
  nand NAND2_1271(II6937,II6939,II6940);
  nand NAND2_1272(II6945,II6921,II6937);
  nand NAND2_1273(II6946,II6921,II6945);
  nand NAND2_1274(II6947,II6937,II6945);
  nand NAND2_1275(WX2223,II6946,II6947);
  nand NAND2_1276(II6954,WX2295,WX2000);
  nand NAND2_1277(II6955,WX2295,II6954);
  nand NAND2_1278(II6956,WX2000,II6954);
  nand NAND2_1279(II6953,II6955,II6956);
  nand NAND2_1280(II6961,WX2064,II6953);
  nand NAND2_1281(II6962,WX2064,II6961);
  nand NAND2_1282(II6963,II6953,II6961);
  nand NAND2_1283(II6952,II6962,II6963);
  nand NAND2_1284(II6969,WX2128,WX2192);
  nand NAND2_1285(II6970,WX2128,II6969);
  nand NAND2_1286(II6971,WX2192,II6969);
  nand NAND2_1287(II6968,II6970,II6971);
  nand NAND2_1288(II6976,II6952,II6968);
  nand NAND2_1289(II6977,II6952,II6976);
  nand NAND2_1290(II6978,II6968,II6976);
  nand NAND2_1291(WX2224,II6977,II6978);
  nand NAND2_1292(II7057,WX1873,WX1778);
  nand NAND2_1293(II7058,WX1873,II7057);
  nand NAND2_1294(II7059,WX1778,II7057);
  nand NAND2_1295(WX2299,II7058,II7059);
  nand NAND2_1296(II7070,WX1874,WX1780);
  nand NAND2_1297(II7071,WX1874,II7070);
  nand NAND2_1298(II7072,WX1780,II7070);
  nand NAND2_1299(WX2306,II7071,II7072);
  nand NAND2_1300(II7083,WX1875,WX1782);
  nand NAND2_1301(II7084,WX1875,II7083);
  nand NAND2_1302(II7085,WX1782,II7083);
  nand NAND2_1303(WX2313,II7084,II7085);
  nand NAND2_1304(II7096,WX1876,WX1784);
  nand NAND2_1305(II7097,WX1876,II7096);
  nand NAND2_1306(II7098,WX1784,II7096);
  nand NAND2_1307(WX2320,II7097,II7098);
  nand NAND2_1308(II7109,WX1877,WX1786);
  nand NAND2_1309(II7110,WX1877,II7109);
  nand NAND2_1310(II7111,WX1786,II7109);
  nand NAND2_1311(WX2327,II7110,II7111);
  nand NAND2_1312(II7122,WX1878,WX1788);
  nand NAND2_1313(II7123,WX1878,II7122);
  nand NAND2_1314(II7124,WX1788,II7122);
  nand NAND2_1315(WX2334,II7123,II7124);
  nand NAND2_1316(II7135,WX1879,WX1790);
  nand NAND2_1317(II7136,WX1879,II7135);
  nand NAND2_1318(II7137,WX1790,II7135);
  nand NAND2_1319(WX2341,II7136,II7137);
  nand NAND2_1320(II7148,WX1880,WX1792);
  nand NAND2_1321(II7149,WX1880,II7148);
  nand NAND2_1322(II7150,WX1792,II7148);
  nand NAND2_1323(WX2348,II7149,II7150);
  nand NAND2_1324(II7161,WX1881,WX1794);
  nand NAND2_1325(II7162,WX1881,II7161);
  nand NAND2_1326(II7163,WX1794,II7161);
  nand NAND2_1327(WX2355,II7162,II7163);
  nand NAND2_1328(II7174,WX1882,WX1796);
  nand NAND2_1329(II7175,WX1882,II7174);
  nand NAND2_1330(II7176,WX1796,II7174);
  nand NAND2_1331(WX2362,II7175,II7176);
  nand NAND2_1332(II7187,WX1883,WX1798);
  nand NAND2_1333(II7188,WX1883,II7187);
  nand NAND2_1334(II7189,WX1798,II7187);
  nand NAND2_1335(WX2369,II7188,II7189);
  nand NAND2_1336(II7200,WX1884,WX1800);
  nand NAND2_1337(II7201,WX1884,II7200);
  nand NAND2_1338(II7202,WX1800,II7200);
  nand NAND2_1339(WX2376,II7201,II7202);
  nand NAND2_1340(II7213,WX1885,WX1802);
  nand NAND2_1341(II7214,WX1885,II7213);
  nand NAND2_1342(II7215,WX1802,II7213);
  nand NAND2_1343(WX2383,II7214,II7215);
  nand NAND2_1344(II7226,WX1886,WX1804);
  nand NAND2_1345(II7227,WX1886,II7226);
  nand NAND2_1346(II7228,WX1804,II7226);
  nand NAND2_1347(WX2390,II7227,II7228);
  nand NAND2_1348(II7239,WX1887,WX1806);
  nand NAND2_1349(II7240,WX1887,II7239);
  nand NAND2_1350(II7241,WX1806,II7239);
  nand NAND2_1351(WX2397,II7240,II7241);
  nand NAND2_1352(II7252,WX1888,WX1808);
  nand NAND2_1353(II7253,WX1888,II7252);
  nand NAND2_1354(II7254,WX1808,II7252);
  nand NAND2_1355(WX2404,II7253,II7254);
  nand NAND2_1356(II7265,WX1889,WX1810);
  nand NAND2_1357(II7266,WX1889,II7265);
  nand NAND2_1358(II7267,WX1810,II7265);
  nand NAND2_1359(WX2411,II7266,II7267);
  nand NAND2_1360(II7278,WX1890,WX1812);
  nand NAND2_1361(II7279,WX1890,II7278);
  nand NAND2_1362(II7280,WX1812,II7278);
  nand NAND2_1363(WX2418,II7279,II7280);
  nand NAND2_1364(II7291,WX1891,WX1814);
  nand NAND2_1365(II7292,WX1891,II7291);
  nand NAND2_1366(II7293,WX1814,II7291);
  nand NAND2_1367(WX2425,II7292,II7293);
  nand NAND2_1368(II7304,WX1892,WX1816);
  nand NAND2_1369(II7305,WX1892,II7304);
  nand NAND2_1370(II7306,WX1816,II7304);
  nand NAND2_1371(WX2432,II7305,II7306);
  nand NAND2_1372(II7317,WX1893,WX1818);
  nand NAND2_1373(II7318,WX1893,II7317);
  nand NAND2_1374(II7319,WX1818,II7317);
  nand NAND2_1375(WX2439,II7318,II7319);
  nand NAND2_1376(II7330,WX1894,WX1820);
  nand NAND2_1377(II7331,WX1894,II7330);
  nand NAND2_1378(II7332,WX1820,II7330);
  nand NAND2_1379(WX2446,II7331,II7332);
  nand NAND2_1380(II7343,WX1895,WX1822);
  nand NAND2_1381(II7344,WX1895,II7343);
  nand NAND2_1382(II7345,WX1822,II7343);
  nand NAND2_1383(WX2453,II7344,II7345);
  nand NAND2_1384(II7356,WX1896,WX1824);
  nand NAND2_1385(II7357,WX1896,II7356);
  nand NAND2_1386(II7358,WX1824,II7356);
  nand NAND2_1387(WX2460,II7357,II7358);
  nand NAND2_1388(II7369,WX1897,WX1826);
  nand NAND2_1389(II7370,WX1897,II7369);
  nand NAND2_1390(II7371,WX1826,II7369);
  nand NAND2_1391(WX2467,II7370,II7371);
  nand NAND2_1392(II7382,WX1898,WX1828);
  nand NAND2_1393(II7383,WX1898,II7382);
  nand NAND2_1394(II7384,WX1828,II7382);
  nand NAND2_1395(WX2474,II7383,II7384);
  nand NAND2_1396(II7395,WX1899,WX1830);
  nand NAND2_1397(II7396,WX1899,II7395);
  nand NAND2_1398(II7397,WX1830,II7395);
  nand NAND2_1399(WX2481,II7396,II7397);
  nand NAND2_1400(II7408,WX1900,WX1832);
  nand NAND2_1401(II7409,WX1900,II7408);
  nand NAND2_1402(II7410,WX1832,II7408);
  nand NAND2_1403(WX2488,II7409,II7410);
  nand NAND2_1404(II7421,WX1901,WX1834);
  nand NAND2_1405(II7422,WX1901,II7421);
  nand NAND2_1406(II7423,WX1834,II7421);
  nand NAND2_1407(WX2495,II7422,II7423);
  nand NAND2_1408(II7434,WX1902,WX1836);
  nand NAND2_1409(II7435,WX1902,II7434);
  nand NAND2_1410(II7436,WX1836,II7434);
  nand NAND2_1411(WX2502,II7435,II7436);
  nand NAND2_1412(II7447,WX1903,WX1838);
  nand NAND2_1413(II7448,WX1903,II7447);
  nand NAND2_1414(II7449,WX1838,II7447);
  nand NAND2_1415(WX2509,II7448,II7449);
  nand NAND2_1416(II7460,WX1904,WX1840);
  nand NAND2_1417(II7461,WX1904,II7460);
  nand NAND2_1418(II7462,WX1840,II7460);
  nand NAND2_1419(WX2516,II7461,II7462);
  nand NAND2_1420(II7475,WX1920,CRC_OUT_8_31);
  nand NAND2_1421(II7476,WX1920,II7475);
  nand NAND2_1422(II7477,CRC_OUT_8_31,II7475);
  nand NAND2_1423(II7474,II7476,II7477);
  nand NAND2_1424(II7482,CRC_OUT_8_15,II7474);
  nand NAND2_1425(II7483,CRC_OUT_8_15,II7482);
  nand NAND2_1426(II7484,II7474,II7482);
  nand NAND2_1427(WX2524,II7483,II7484);
  nand NAND2_1428(II7490,WX1925,CRC_OUT_8_31);
  nand NAND2_1429(II7491,WX1925,II7490);
  nand NAND2_1430(II7492,CRC_OUT_8_31,II7490);
  nand NAND2_1431(II7489,II7491,II7492);
  nand NAND2_1432(II7497,CRC_OUT_8_10,II7489);
  nand NAND2_1433(II7498,CRC_OUT_8_10,II7497);
  nand NAND2_1434(II7499,II7489,II7497);
  nand NAND2_1435(WX2525,II7498,II7499);
  nand NAND2_1436(II7505,WX1932,CRC_OUT_8_31);
  nand NAND2_1437(II7506,WX1932,II7505);
  nand NAND2_1438(II7507,CRC_OUT_8_31,II7505);
  nand NAND2_1439(II7504,II7506,II7507);
  nand NAND2_1440(II7512,CRC_OUT_8_3,II7504);
  nand NAND2_1441(II7513,CRC_OUT_8_3,II7512);
  nand NAND2_1442(II7514,II7504,II7512);
  nand NAND2_1443(WX2526,II7513,II7514);
  nand NAND2_1444(II7519,WX1936,CRC_OUT_8_31);
  nand NAND2_1445(II7520,WX1936,II7519);
  nand NAND2_1446(II7521,CRC_OUT_8_31,II7519);
  nand NAND2_1447(WX2527,II7520,II7521);
  nand NAND2_1448(II7526,WX1905,CRC_OUT_8_30);
  nand NAND2_1449(II7527,WX1905,II7526);
  nand NAND2_1450(II7528,CRC_OUT_8_30,II7526);
  nand NAND2_1451(WX2528,II7527,II7528);
  nand NAND2_1452(II7533,WX1906,CRC_OUT_8_29);
  nand NAND2_1453(II7534,WX1906,II7533);
  nand NAND2_1454(II7535,CRC_OUT_8_29,II7533);
  nand NAND2_1455(WX2529,II7534,II7535);
  nand NAND2_1456(II7540,WX1907,CRC_OUT_8_28);
  nand NAND2_1457(II7541,WX1907,II7540);
  nand NAND2_1458(II7542,CRC_OUT_8_28,II7540);
  nand NAND2_1459(WX2530,II7541,II7542);
  nand NAND2_1460(II7547,WX1908,CRC_OUT_8_27);
  nand NAND2_1461(II7548,WX1908,II7547);
  nand NAND2_1462(II7549,CRC_OUT_8_27,II7547);
  nand NAND2_1463(WX2531,II7548,II7549);
  nand NAND2_1464(II7554,WX1909,CRC_OUT_8_26);
  nand NAND2_1465(II7555,WX1909,II7554);
  nand NAND2_1466(II7556,CRC_OUT_8_26,II7554);
  nand NAND2_1467(WX2532,II7555,II7556);
  nand NAND2_1468(II7561,WX1910,CRC_OUT_8_25);
  nand NAND2_1469(II7562,WX1910,II7561);
  nand NAND2_1470(II7563,CRC_OUT_8_25,II7561);
  nand NAND2_1471(WX2533,II7562,II7563);
  nand NAND2_1472(II7568,WX1911,CRC_OUT_8_24);
  nand NAND2_1473(II7569,WX1911,II7568);
  nand NAND2_1474(II7570,CRC_OUT_8_24,II7568);
  nand NAND2_1475(WX2534,II7569,II7570);
  nand NAND2_1476(II7575,WX1912,CRC_OUT_8_23);
  nand NAND2_1477(II7576,WX1912,II7575);
  nand NAND2_1478(II7577,CRC_OUT_8_23,II7575);
  nand NAND2_1479(WX2535,II7576,II7577);
  nand NAND2_1480(II7582,WX1913,CRC_OUT_8_22);
  nand NAND2_1481(II7583,WX1913,II7582);
  nand NAND2_1482(II7584,CRC_OUT_8_22,II7582);
  nand NAND2_1483(WX2536,II7583,II7584);
  nand NAND2_1484(II7589,WX1914,CRC_OUT_8_21);
  nand NAND2_1485(II7590,WX1914,II7589);
  nand NAND2_1486(II7591,CRC_OUT_8_21,II7589);
  nand NAND2_1487(WX2537,II7590,II7591);
  nand NAND2_1488(II7596,WX1915,CRC_OUT_8_20);
  nand NAND2_1489(II7597,WX1915,II7596);
  nand NAND2_1490(II7598,CRC_OUT_8_20,II7596);
  nand NAND2_1491(WX2538,II7597,II7598);
  nand NAND2_1492(II7603,WX1916,CRC_OUT_8_19);
  nand NAND2_1493(II7604,WX1916,II7603);
  nand NAND2_1494(II7605,CRC_OUT_8_19,II7603);
  nand NAND2_1495(WX2539,II7604,II7605);
  nand NAND2_1496(II7610,WX1917,CRC_OUT_8_18);
  nand NAND2_1497(II7611,WX1917,II7610);
  nand NAND2_1498(II7612,CRC_OUT_8_18,II7610);
  nand NAND2_1499(WX2540,II7611,II7612);
  nand NAND2_1500(II7617,WX1918,CRC_OUT_8_17);
  nand NAND2_1501(II7618,WX1918,II7617);
  nand NAND2_1502(II7619,CRC_OUT_8_17,II7617);
  nand NAND2_1503(WX2541,II7618,II7619);
  nand NAND2_1504(II7624,WX1919,CRC_OUT_8_16);
  nand NAND2_1505(II7625,WX1919,II7624);
  nand NAND2_1506(II7626,CRC_OUT_8_16,II7624);
  nand NAND2_1507(WX2542,II7625,II7626);
  nand NAND2_1508(II7631,WX1921,CRC_OUT_8_14);
  nand NAND2_1509(II7632,WX1921,II7631);
  nand NAND2_1510(II7633,CRC_OUT_8_14,II7631);
  nand NAND2_1511(WX2543,II7632,II7633);
  nand NAND2_1512(II7638,WX1922,CRC_OUT_8_13);
  nand NAND2_1513(II7639,WX1922,II7638);
  nand NAND2_1514(II7640,CRC_OUT_8_13,II7638);
  nand NAND2_1515(WX2544,II7639,II7640);
  nand NAND2_1516(II7645,WX1923,CRC_OUT_8_12);
  nand NAND2_1517(II7646,WX1923,II7645);
  nand NAND2_1518(II7647,CRC_OUT_8_12,II7645);
  nand NAND2_1519(WX2545,II7646,II7647);
  nand NAND2_1520(II7652,WX1924,CRC_OUT_8_11);
  nand NAND2_1521(II7653,WX1924,II7652);
  nand NAND2_1522(II7654,CRC_OUT_8_11,II7652);
  nand NAND2_1523(WX2546,II7653,II7654);
  nand NAND2_1524(II7659,WX1926,CRC_OUT_8_9);
  nand NAND2_1525(II7660,WX1926,II7659);
  nand NAND2_1526(II7661,CRC_OUT_8_9,II7659);
  nand NAND2_1527(WX2547,II7660,II7661);
  nand NAND2_1528(II7666,WX1927,CRC_OUT_8_8);
  nand NAND2_1529(II7667,WX1927,II7666);
  nand NAND2_1530(II7668,CRC_OUT_8_8,II7666);
  nand NAND2_1531(WX2548,II7667,II7668);
  nand NAND2_1532(II7673,WX1928,CRC_OUT_8_7);
  nand NAND2_1533(II7674,WX1928,II7673);
  nand NAND2_1534(II7675,CRC_OUT_8_7,II7673);
  nand NAND2_1535(WX2549,II7674,II7675);
  nand NAND2_1536(II7680,WX1929,CRC_OUT_8_6);
  nand NAND2_1537(II7681,WX1929,II7680);
  nand NAND2_1538(II7682,CRC_OUT_8_6,II7680);
  nand NAND2_1539(WX2550,II7681,II7682);
  nand NAND2_1540(II7687,WX1930,CRC_OUT_8_5);
  nand NAND2_1541(II7688,WX1930,II7687);
  nand NAND2_1542(II7689,CRC_OUT_8_5,II7687);
  nand NAND2_1543(WX2551,II7688,II7689);
  nand NAND2_1544(II7694,WX1931,CRC_OUT_8_4);
  nand NAND2_1545(II7695,WX1931,II7694);
  nand NAND2_1546(II7696,CRC_OUT_8_4,II7694);
  nand NAND2_1547(WX2552,II7695,II7696);
  nand NAND2_1548(II7701,WX1933,CRC_OUT_8_2);
  nand NAND2_1549(II7702,WX1933,II7701);
  nand NAND2_1550(II7703,CRC_OUT_8_2,II7701);
  nand NAND2_1551(WX2553,II7702,II7703);
  nand NAND2_1552(II7708,WX1934,CRC_OUT_8_1);
  nand NAND2_1553(II7709,WX1934,II7708);
  nand NAND2_1554(II7710,CRC_OUT_8_1,II7708);
  nand NAND2_1555(WX2554,II7709,II7710);
  nand NAND2_1556(II7715,WX1935,CRC_OUT_8_0);
  nand NAND2_1557(II7716,WX1935,II7715);
  nand NAND2_1558(II7717,CRC_OUT_8_0,II7715);
  nand NAND2_1559(WX2555,II7716,II7717);
  nand NAND2_1560(II9998,WX3587,WX3231);
  nand NAND2_1561(II9999,WX3587,II9998);
  nand NAND2_1562(II10000,WX3231,II9998);
  nand NAND2_1563(II9997,II9999,II10000);
  nand NAND2_1564(II10005,WX3295,II9997);
  nand NAND2_1565(II10006,WX3295,II10005);
  nand NAND2_1566(II10007,II9997,II10005);
  nand NAND2_1567(II9996,II10006,II10007);
  nand NAND2_1568(II10013,WX3359,WX3423);
  nand NAND2_1569(II10014,WX3359,II10013);
  nand NAND2_1570(II10015,WX3423,II10013);
  nand NAND2_1571(II10012,II10014,II10015);
  nand NAND2_1572(II10020,II9996,II10012);
  nand NAND2_1573(II10021,II9996,II10020);
  nand NAND2_1574(II10022,II10012,II10020);
  nand NAND2_1575(WX3486,II10021,II10022);
  nand NAND2_1576(II10029,WX3587,WX3233);
  nand NAND2_1577(II10030,WX3587,II10029);
  nand NAND2_1578(II10031,WX3233,II10029);
  nand NAND2_1579(II10028,II10030,II10031);
  nand NAND2_1580(II10036,WX3297,II10028);
  nand NAND2_1581(II10037,WX3297,II10036);
  nand NAND2_1582(II10038,II10028,II10036);
  nand NAND2_1583(II10027,II10037,II10038);
  nand NAND2_1584(II10044,WX3361,WX3425);
  nand NAND2_1585(II10045,WX3361,II10044);
  nand NAND2_1586(II10046,WX3425,II10044);
  nand NAND2_1587(II10043,II10045,II10046);
  nand NAND2_1588(II10051,II10027,II10043);
  nand NAND2_1589(II10052,II10027,II10051);
  nand NAND2_1590(II10053,II10043,II10051);
  nand NAND2_1591(WX3487,II10052,II10053);
  nand NAND2_1592(II10060,WX3587,WX3235);
  nand NAND2_1593(II10061,WX3587,II10060);
  nand NAND2_1594(II10062,WX3235,II10060);
  nand NAND2_1595(II10059,II10061,II10062);
  nand NAND2_1596(II10067,WX3299,II10059);
  nand NAND2_1597(II10068,WX3299,II10067);
  nand NAND2_1598(II10069,II10059,II10067);
  nand NAND2_1599(II10058,II10068,II10069);
  nand NAND2_1600(II10075,WX3363,WX3427);
  nand NAND2_1601(II10076,WX3363,II10075);
  nand NAND2_1602(II10077,WX3427,II10075);
  nand NAND2_1603(II10074,II10076,II10077);
  nand NAND2_1604(II10082,II10058,II10074);
  nand NAND2_1605(II10083,II10058,II10082);
  nand NAND2_1606(II10084,II10074,II10082);
  nand NAND2_1607(WX3488,II10083,II10084);
  nand NAND2_1608(II10091,WX3587,WX3237);
  nand NAND2_1609(II10092,WX3587,II10091);
  nand NAND2_1610(II10093,WX3237,II10091);
  nand NAND2_1611(II10090,II10092,II10093);
  nand NAND2_1612(II10098,WX3301,II10090);
  nand NAND2_1613(II10099,WX3301,II10098);
  nand NAND2_1614(II10100,II10090,II10098);
  nand NAND2_1615(II10089,II10099,II10100);
  nand NAND2_1616(II10106,WX3365,WX3429);
  nand NAND2_1617(II10107,WX3365,II10106);
  nand NAND2_1618(II10108,WX3429,II10106);
  nand NAND2_1619(II10105,II10107,II10108);
  nand NAND2_1620(II10113,II10089,II10105);
  nand NAND2_1621(II10114,II10089,II10113);
  nand NAND2_1622(II10115,II10105,II10113);
  nand NAND2_1623(WX3489,II10114,II10115);
  nand NAND2_1624(II10122,WX3587,WX3239);
  nand NAND2_1625(II10123,WX3587,II10122);
  nand NAND2_1626(II10124,WX3239,II10122);
  nand NAND2_1627(II10121,II10123,II10124);
  nand NAND2_1628(II10129,WX3303,II10121);
  nand NAND2_1629(II10130,WX3303,II10129);
  nand NAND2_1630(II10131,II10121,II10129);
  nand NAND2_1631(II10120,II10130,II10131);
  nand NAND2_1632(II10137,WX3367,WX3431);
  nand NAND2_1633(II10138,WX3367,II10137);
  nand NAND2_1634(II10139,WX3431,II10137);
  nand NAND2_1635(II10136,II10138,II10139);
  nand NAND2_1636(II10144,II10120,II10136);
  nand NAND2_1637(II10145,II10120,II10144);
  nand NAND2_1638(II10146,II10136,II10144);
  nand NAND2_1639(WX3490,II10145,II10146);
  nand NAND2_1640(II10153,WX3587,WX3241);
  nand NAND2_1641(II10154,WX3587,II10153);
  nand NAND2_1642(II10155,WX3241,II10153);
  nand NAND2_1643(II10152,II10154,II10155);
  nand NAND2_1644(II10160,WX3305,II10152);
  nand NAND2_1645(II10161,WX3305,II10160);
  nand NAND2_1646(II10162,II10152,II10160);
  nand NAND2_1647(II10151,II10161,II10162);
  nand NAND2_1648(II10168,WX3369,WX3433);
  nand NAND2_1649(II10169,WX3369,II10168);
  nand NAND2_1650(II10170,WX3433,II10168);
  nand NAND2_1651(II10167,II10169,II10170);
  nand NAND2_1652(II10175,II10151,II10167);
  nand NAND2_1653(II10176,II10151,II10175);
  nand NAND2_1654(II10177,II10167,II10175);
  nand NAND2_1655(WX3491,II10176,II10177);
  nand NAND2_1656(II10184,WX3587,WX3243);
  nand NAND2_1657(II10185,WX3587,II10184);
  nand NAND2_1658(II10186,WX3243,II10184);
  nand NAND2_1659(II10183,II10185,II10186);
  nand NAND2_1660(II10191,WX3307,II10183);
  nand NAND2_1661(II10192,WX3307,II10191);
  nand NAND2_1662(II10193,II10183,II10191);
  nand NAND2_1663(II10182,II10192,II10193);
  nand NAND2_1664(II10199,WX3371,WX3435);
  nand NAND2_1665(II10200,WX3371,II10199);
  nand NAND2_1666(II10201,WX3435,II10199);
  nand NAND2_1667(II10198,II10200,II10201);
  nand NAND2_1668(II10206,II10182,II10198);
  nand NAND2_1669(II10207,II10182,II10206);
  nand NAND2_1670(II10208,II10198,II10206);
  nand NAND2_1671(WX3492,II10207,II10208);
  nand NAND2_1672(II10215,WX3587,WX3245);
  nand NAND2_1673(II10216,WX3587,II10215);
  nand NAND2_1674(II10217,WX3245,II10215);
  nand NAND2_1675(II10214,II10216,II10217);
  nand NAND2_1676(II10222,WX3309,II10214);
  nand NAND2_1677(II10223,WX3309,II10222);
  nand NAND2_1678(II10224,II10214,II10222);
  nand NAND2_1679(II10213,II10223,II10224);
  nand NAND2_1680(II10230,WX3373,WX3437);
  nand NAND2_1681(II10231,WX3373,II10230);
  nand NAND2_1682(II10232,WX3437,II10230);
  nand NAND2_1683(II10229,II10231,II10232);
  nand NAND2_1684(II10237,II10213,II10229);
  nand NAND2_1685(II10238,II10213,II10237);
  nand NAND2_1686(II10239,II10229,II10237);
  nand NAND2_1687(WX3493,II10238,II10239);
  nand NAND2_1688(II10246,WX3587,WX3247);
  nand NAND2_1689(II10247,WX3587,II10246);
  nand NAND2_1690(II10248,WX3247,II10246);
  nand NAND2_1691(II10245,II10247,II10248);
  nand NAND2_1692(II10253,WX3311,II10245);
  nand NAND2_1693(II10254,WX3311,II10253);
  nand NAND2_1694(II10255,II10245,II10253);
  nand NAND2_1695(II10244,II10254,II10255);
  nand NAND2_1696(II10261,WX3375,WX3439);
  nand NAND2_1697(II10262,WX3375,II10261);
  nand NAND2_1698(II10263,WX3439,II10261);
  nand NAND2_1699(II10260,II10262,II10263);
  nand NAND2_1700(II10268,II10244,II10260);
  nand NAND2_1701(II10269,II10244,II10268);
  nand NAND2_1702(II10270,II10260,II10268);
  nand NAND2_1703(WX3494,II10269,II10270);
  nand NAND2_1704(II10277,WX3587,WX3249);
  nand NAND2_1705(II10278,WX3587,II10277);
  nand NAND2_1706(II10279,WX3249,II10277);
  nand NAND2_1707(II10276,II10278,II10279);
  nand NAND2_1708(II10284,WX3313,II10276);
  nand NAND2_1709(II10285,WX3313,II10284);
  nand NAND2_1710(II10286,II10276,II10284);
  nand NAND2_1711(II10275,II10285,II10286);
  nand NAND2_1712(II10292,WX3377,WX3441);
  nand NAND2_1713(II10293,WX3377,II10292);
  nand NAND2_1714(II10294,WX3441,II10292);
  nand NAND2_1715(II10291,II10293,II10294);
  nand NAND2_1716(II10299,II10275,II10291);
  nand NAND2_1717(II10300,II10275,II10299);
  nand NAND2_1718(II10301,II10291,II10299);
  nand NAND2_1719(WX3495,II10300,II10301);
  nand NAND2_1720(II10308,WX3587,WX3251);
  nand NAND2_1721(II10309,WX3587,II10308);
  nand NAND2_1722(II10310,WX3251,II10308);
  nand NAND2_1723(II10307,II10309,II10310);
  nand NAND2_1724(II10315,WX3315,II10307);
  nand NAND2_1725(II10316,WX3315,II10315);
  nand NAND2_1726(II10317,II10307,II10315);
  nand NAND2_1727(II10306,II10316,II10317);
  nand NAND2_1728(II10323,WX3379,WX3443);
  nand NAND2_1729(II10324,WX3379,II10323);
  nand NAND2_1730(II10325,WX3443,II10323);
  nand NAND2_1731(II10322,II10324,II10325);
  nand NAND2_1732(II10330,II10306,II10322);
  nand NAND2_1733(II10331,II10306,II10330);
  nand NAND2_1734(II10332,II10322,II10330);
  nand NAND2_1735(WX3496,II10331,II10332);
  nand NAND2_1736(II10339,WX3587,WX3253);
  nand NAND2_1737(II10340,WX3587,II10339);
  nand NAND2_1738(II10341,WX3253,II10339);
  nand NAND2_1739(II10338,II10340,II10341);
  nand NAND2_1740(II10346,WX3317,II10338);
  nand NAND2_1741(II10347,WX3317,II10346);
  nand NAND2_1742(II10348,II10338,II10346);
  nand NAND2_1743(II10337,II10347,II10348);
  nand NAND2_1744(II10354,WX3381,WX3445);
  nand NAND2_1745(II10355,WX3381,II10354);
  nand NAND2_1746(II10356,WX3445,II10354);
  nand NAND2_1747(II10353,II10355,II10356);
  nand NAND2_1748(II10361,II10337,II10353);
  nand NAND2_1749(II10362,II10337,II10361);
  nand NAND2_1750(II10363,II10353,II10361);
  nand NAND2_1751(WX3497,II10362,II10363);
  nand NAND2_1752(II10370,WX3587,WX3255);
  nand NAND2_1753(II10371,WX3587,II10370);
  nand NAND2_1754(II10372,WX3255,II10370);
  nand NAND2_1755(II10369,II10371,II10372);
  nand NAND2_1756(II10377,WX3319,II10369);
  nand NAND2_1757(II10378,WX3319,II10377);
  nand NAND2_1758(II10379,II10369,II10377);
  nand NAND2_1759(II10368,II10378,II10379);
  nand NAND2_1760(II10385,WX3383,WX3447);
  nand NAND2_1761(II10386,WX3383,II10385);
  nand NAND2_1762(II10387,WX3447,II10385);
  nand NAND2_1763(II10384,II10386,II10387);
  nand NAND2_1764(II10392,II10368,II10384);
  nand NAND2_1765(II10393,II10368,II10392);
  nand NAND2_1766(II10394,II10384,II10392);
  nand NAND2_1767(WX3498,II10393,II10394);
  nand NAND2_1768(II10401,WX3587,WX3257);
  nand NAND2_1769(II10402,WX3587,II10401);
  nand NAND2_1770(II10403,WX3257,II10401);
  nand NAND2_1771(II10400,II10402,II10403);
  nand NAND2_1772(II10408,WX3321,II10400);
  nand NAND2_1773(II10409,WX3321,II10408);
  nand NAND2_1774(II10410,II10400,II10408);
  nand NAND2_1775(II10399,II10409,II10410);
  nand NAND2_1776(II10416,WX3385,WX3449);
  nand NAND2_1777(II10417,WX3385,II10416);
  nand NAND2_1778(II10418,WX3449,II10416);
  nand NAND2_1779(II10415,II10417,II10418);
  nand NAND2_1780(II10423,II10399,II10415);
  nand NAND2_1781(II10424,II10399,II10423);
  nand NAND2_1782(II10425,II10415,II10423);
  nand NAND2_1783(WX3499,II10424,II10425);
  nand NAND2_1784(II10432,WX3587,WX3259);
  nand NAND2_1785(II10433,WX3587,II10432);
  nand NAND2_1786(II10434,WX3259,II10432);
  nand NAND2_1787(II10431,II10433,II10434);
  nand NAND2_1788(II10439,WX3323,II10431);
  nand NAND2_1789(II10440,WX3323,II10439);
  nand NAND2_1790(II10441,II10431,II10439);
  nand NAND2_1791(II10430,II10440,II10441);
  nand NAND2_1792(II10447,WX3387,WX3451);
  nand NAND2_1793(II10448,WX3387,II10447);
  nand NAND2_1794(II10449,WX3451,II10447);
  nand NAND2_1795(II10446,II10448,II10449);
  nand NAND2_1796(II10454,II10430,II10446);
  nand NAND2_1797(II10455,II10430,II10454);
  nand NAND2_1798(II10456,II10446,II10454);
  nand NAND2_1799(WX3500,II10455,II10456);
  nand NAND2_1800(II10463,WX3587,WX3261);
  nand NAND2_1801(II10464,WX3587,II10463);
  nand NAND2_1802(II10465,WX3261,II10463);
  nand NAND2_1803(II10462,II10464,II10465);
  nand NAND2_1804(II10470,WX3325,II10462);
  nand NAND2_1805(II10471,WX3325,II10470);
  nand NAND2_1806(II10472,II10462,II10470);
  nand NAND2_1807(II10461,II10471,II10472);
  nand NAND2_1808(II10478,WX3389,WX3453);
  nand NAND2_1809(II10479,WX3389,II10478);
  nand NAND2_1810(II10480,WX3453,II10478);
  nand NAND2_1811(II10477,II10479,II10480);
  nand NAND2_1812(II10485,II10461,II10477);
  nand NAND2_1813(II10486,II10461,II10485);
  nand NAND2_1814(II10487,II10477,II10485);
  nand NAND2_1815(WX3501,II10486,II10487);
  nand NAND2_1816(II10494,WX3588,WX3263);
  nand NAND2_1817(II10495,WX3588,II10494);
  nand NAND2_1818(II10496,WX3263,II10494);
  nand NAND2_1819(II10493,II10495,II10496);
  nand NAND2_1820(II10501,WX3327,II10493);
  nand NAND2_1821(II10502,WX3327,II10501);
  nand NAND2_1822(II10503,II10493,II10501);
  nand NAND2_1823(II10492,II10502,II10503);
  nand NAND2_1824(II10509,WX3391,WX3455);
  nand NAND2_1825(II10510,WX3391,II10509);
  nand NAND2_1826(II10511,WX3455,II10509);
  nand NAND2_1827(II10508,II10510,II10511);
  nand NAND2_1828(II10516,II10492,II10508);
  nand NAND2_1829(II10517,II10492,II10516);
  nand NAND2_1830(II10518,II10508,II10516);
  nand NAND2_1831(WX3502,II10517,II10518);
  nand NAND2_1832(II10525,WX3588,WX3265);
  nand NAND2_1833(II10526,WX3588,II10525);
  nand NAND2_1834(II10527,WX3265,II10525);
  nand NAND2_1835(II10524,II10526,II10527);
  nand NAND2_1836(II10532,WX3329,II10524);
  nand NAND2_1837(II10533,WX3329,II10532);
  nand NAND2_1838(II10534,II10524,II10532);
  nand NAND2_1839(II10523,II10533,II10534);
  nand NAND2_1840(II10540,WX3393,WX3457);
  nand NAND2_1841(II10541,WX3393,II10540);
  nand NAND2_1842(II10542,WX3457,II10540);
  nand NAND2_1843(II10539,II10541,II10542);
  nand NAND2_1844(II10547,II10523,II10539);
  nand NAND2_1845(II10548,II10523,II10547);
  nand NAND2_1846(II10549,II10539,II10547);
  nand NAND2_1847(WX3503,II10548,II10549);
  nand NAND2_1848(II10556,WX3588,WX3267);
  nand NAND2_1849(II10557,WX3588,II10556);
  nand NAND2_1850(II10558,WX3267,II10556);
  nand NAND2_1851(II10555,II10557,II10558);
  nand NAND2_1852(II10563,WX3331,II10555);
  nand NAND2_1853(II10564,WX3331,II10563);
  nand NAND2_1854(II10565,II10555,II10563);
  nand NAND2_1855(II10554,II10564,II10565);
  nand NAND2_1856(II10571,WX3395,WX3459);
  nand NAND2_1857(II10572,WX3395,II10571);
  nand NAND2_1858(II10573,WX3459,II10571);
  nand NAND2_1859(II10570,II10572,II10573);
  nand NAND2_1860(II10578,II10554,II10570);
  nand NAND2_1861(II10579,II10554,II10578);
  nand NAND2_1862(II10580,II10570,II10578);
  nand NAND2_1863(WX3504,II10579,II10580);
  nand NAND2_1864(II10587,WX3588,WX3269);
  nand NAND2_1865(II10588,WX3588,II10587);
  nand NAND2_1866(II10589,WX3269,II10587);
  nand NAND2_1867(II10586,II10588,II10589);
  nand NAND2_1868(II10594,WX3333,II10586);
  nand NAND2_1869(II10595,WX3333,II10594);
  nand NAND2_1870(II10596,II10586,II10594);
  nand NAND2_1871(II10585,II10595,II10596);
  nand NAND2_1872(II10602,WX3397,WX3461);
  nand NAND2_1873(II10603,WX3397,II10602);
  nand NAND2_1874(II10604,WX3461,II10602);
  nand NAND2_1875(II10601,II10603,II10604);
  nand NAND2_1876(II10609,II10585,II10601);
  nand NAND2_1877(II10610,II10585,II10609);
  nand NAND2_1878(II10611,II10601,II10609);
  nand NAND2_1879(WX3505,II10610,II10611);
  nand NAND2_1880(II10618,WX3588,WX3271);
  nand NAND2_1881(II10619,WX3588,II10618);
  nand NAND2_1882(II10620,WX3271,II10618);
  nand NAND2_1883(II10617,II10619,II10620);
  nand NAND2_1884(II10625,WX3335,II10617);
  nand NAND2_1885(II10626,WX3335,II10625);
  nand NAND2_1886(II10627,II10617,II10625);
  nand NAND2_1887(II10616,II10626,II10627);
  nand NAND2_1888(II10633,WX3399,WX3463);
  nand NAND2_1889(II10634,WX3399,II10633);
  nand NAND2_1890(II10635,WX3463,II10633);
  nand NAND2_1891(II10632,II10634,II10635);
  nand NAND2_1892(II10640,II10616,II10632);
  nand NAND2_1893(II10641,II10616,II10640);
  nand NAND2_1894(II10642,II10632,II10640);
  nand NAND2_1895(WX3506,II10641,II10642);
  nand NAND2_1896(II10649,WX3588,WX3273);
  nand NAND2_1897(II10650,WX3588,II10649);
  nand NAND2_1898(II10651,WX3273,II10649);
  nand NAND2_1899(II10648,II10650,II10651);
  nand NAND2_1900(II10656,WX3337,II10648);
  nand NAND2_1901(II10657,WX3337,II10656);
  nand NAND2_1902(II10658,II10648,II10656);
  nand NAND2_1903(II10647,II10657,II10658);
  nand NAND2_1904(II10664,WX3401,WX3465);
  nand NAND2_1905(II10665,WX3401,II10664);
  nand NAND2_1906(II10666,WX3465,II10664);
  nand NAND2_1907(II10663,II10665,II10666);
  nand NAND2_1908(II10671,II10647,II10663);
  nand NAND2_1909(II10672,II10647,II10671);
  nand NAND2_1910(II10673,II10663,II10671);
  nand NAND2_1911(WX3507,II10672,II10673);
  nand NAND2_1912(II10680,WX3588,WX3275);
  nand NAND2_1913(II10681,WX3588,II10680);
  nand NAND2_1914(II10682,WX3275,II10680);
  nand NAND2_1915(II10679,II10681,II10682);
  nand NAND2_1916(II10687,WX3339,II10679);
  nand NAND2_1917(II10688,WX3339,II10687);
  nand NAND2_1918(II10689,II10679,II10687);
  nand NAND2_1919(II10678,II10688,II10689);
  nand NAND2_1920(II10695,WX3403,WX3467);
  nand NAND2_1921(II10696,WX3403,II10695);
  nand NAND2_1922(II10697,WX3467,II10695);
  nand NAND2_1923(II10694,II10696,II10697);
  nand NAND2_1924(II10702,II10678,II10694);
  nand NAND2_1925(II10703,II10678,II10702);
  nand NAND2_1926(II10704,II10694,II10702);
  nand NAND2_1927(WX3508,II10703,II10704);
  nand NAND2_1928(II10711,WX3588,WX3277);
  nand NAND2_1929(II10712,WX3588,II10711);
  nand NAND2_1930(II10713,WX3277,II10711);
  nand NAND2_1931(II10710,II10712,II10713);
  nand NAND2_1932(II10718,WX3341,II10710);
  nand NAND2_1933(II10719,WX3341,II10718);
  nand NAND2_1934(II10720,II10710,II10718);
  nand NAND2_1935(II10709,II10719,II10720);
  nand NAND2_1936(II10726,WX3405,WX3469);
  nand NAND2_1937(II10727,WX3405,II10726);
  nand NAND2_1938(II10728,WX3469,II10726);
  nand NAND2_1939(II10725,II10727,II10728);
  nand NAND2_1940(II10733,II10709,II10725);
  nand NAND2_1941(II10734,II10709,II10733);
  nand NAND2_1942(II10735,II10725,II10733);
  nand NAND2_1943(WX3509,II10734,II10735);
  nand NAND2_1944(II10742,WX3588,WX3279);
  nand NAND2_1945(II10743,WX3588,II10742);
  nand NAND2_1946(II10744,WX3279,II10742);
  nand NAND2_1947(II10741,II10743,II10744);
  nand NAND2_1948(II10749,WX3343,II10741);
  nand NAND2_1949(II10750,WX3343,II10749);
  nand NAND2_1950(II10751,II10741,II10749);
  nand NAND2_1951(II10740,II10750,II10751);
  nand NAND2_1952(II10757,WX3407,WX3471);
  nand NAND2_1953(II10758,WX3407,II10757);
  nand NAND2_1954(II10759,WX3471,II10757);
  nand NAND2_1955(II10756,II10758,II10759);
  nand NAND2_1956(II10764,II10740,II10756);
  nand NAND2_1957(II10765,II10740,II10764);
  nand NAND2_1958(II10766,II10756,II10764);
  nand NAND2_1959(WX3510,II10765,II10766);
  nand NAND2_1960(II10773,WX3588,WX3281);
  nand NAND2_1961(II10774,WX3588,II10773);
  nand NAND2_1962(II10775,WX3281,II10773);
  nand NAND2_1963(II10772,II10774,II10775);
  nand NAND2_1964(II10780,WX3345,II10772);
  nand NAND2_1965(II10781,WX3345,II10780);
  nand NAND2_1966(II10782,II10772,II10780);
  nand NAND2_1967(II10771,II10781,II10782);
  nand NAND2_1968(II10788,WX3409,WX3473);
  nand NAND2_1969(II10789,WX3409,II10788);
  nand NAND2_1970(II10790,WX3473,II10788);
  nand NAND2_1971(II10787,II10789,II10790);
  nand NAND2_1972(II10795,II10771,II10787);
  nand NAND2_1973(II10796,II10771,II10795);
  nand NAND2_1974(II10797,II10787,II10795);
  nand NAND2_1975(WX3511,II10796,II10797);
  nand NAND2_1976(II10804,WX3588,WX3283);
  nand NAND2_1977(II10805,WX3588,II10804);
  nand NAND2_1978(II10806,WX3283,II10804);
  nand NAND2_1979(II10803,II10805,II10806);
  nand NAND2_1980(II10811,WX3347,II10803);
  nand NAND2_1981(II10812,WX3347,II10811);
  nand NAND2_1982(II10813,II10803,II10811);
  nand NAND2_1983(II10802,II10812,II10813);
  nand NAND2_1984(II10819,WX3411,WX3475);
  nand NAND2_1985(II10820,WX3411,II10819);
  nand NAND2_1986(II10821,WX3475,II10819);
  nand NAND2_1987(II10818,II10820,II10821);
  nand NAND2_1988(II10826,II10802,II10818);
  nand NAND2_1989(II10827,II10802,II10826);
  nand NAND2_1990(II10828,II10818,II10826);
  nand NAND2_1991(WX3512,II10827,II10828);
  nand NAND2_1992(II10835,WX3588,WX3285);
  nand NAND2_1993(II10836,WX3588,II10835);
  nand NAND2_1994(II10837,WX3285,II10835);
  nand NAND2_1995(II10834,II10836,II10837);
  nand NAND2_1996(II10842,WX3349,II10834);
  nand NAND2_1997(II10843,WX3349,II10842);
  nand NAND2_1998(II10844,II10834,II10842);
  nand NAND2_1999(II10833,II10843,II10844);
  nand NAND2_2000(II10850,WX3413,WX3477);
  nand NAND2_2001(II10851,WX3413,II10850);
  nand NAND2_2002(II10852,WX3477,II10850);
  nand NAND2_2003(II10849,II10851,II10852);
  nand NAND2_2004(II10857,II10833,II10849);
  nand NAND2_2005(II10858,II10833,II10857);
  nand NAND2_2006(II10859,II10849,II10857);
  nand NAND2_2007(WX3513,II10858,II10859);
  nand NAND2_2008(II10866,WX3588,WX3287);
  nand NAND2_2009(II10867,WX3588,II10866);
  nand NAND2_2010(II10868,WX3287,II10866);
  nand NAND2_2011(II10865,II10867,II10868);
  nand NAND2_2012(II10873,WX3351,II10865);
  nand NAND2_2013(II10874,WX3351,II10873);
  nand NAND2_2014(II10875,II10865,II10873);
  nand NAND2_2015(II10864,II10874,II10875);
  nand NAND2_2016(II10881,WX3415,WX3479);
  nand NAND2_2017(II10882,WX3415,II10881);
  nand NAND2_2018(II10883,WX3479,II10881);
  nand NAND2_2019(II10880,II10882,II10883);
  nand NAND2_2020(II10888,II10864,II10880);
  nand NAND2_2021(II10889,II10864,II10888);
  nand NAND2_2022(II10890,II10880,II10888);
  nand NAND2_2023(WX3514,II10889,II10890);
  nand NAND2_2024(II10897,WX3588,WX3289);
  nand NAND2_2025(II10898,WX3588,II10897);
  nand NAND2_2026(II10899,WX3289,II10897);
  nand NAND2_2027(II10896,II10898,II10899);
  nand NAND2_2028(II10904,WX3353,II10896);
  nand NAND2_2029(II10905,WX3353,II10904);
  nand NAND2_2030(II10906,II10896,II10904);
  nand NAND2_2031(II10895,II10905,II10906);
  nand NAND2_2032(II10912,WX3417,WX3481);
  nand NAND2_2033(II10913,WX3417,II10912);
  nand NAND2_2034(II10914,WX3481,II10912);
  nand NAND2_2035(II10911,II10913,II10914);
  nand NAND2_2036(II10919,II10895,II10911);
  nand NAND2_2037(II10920,II10895,II10919);
  nand NAND2_2038(II10921,II10911,II10919);
  nand NAND2_2039(WX3515,II10920,II10921);
  nand NAND2_2040(II10928,WX3588,WX3291);
  nand NAND2_2041(II10929,WX3588,II10928);
  nand NAND2_2042(II10930,WX3291,II10928);
  nand NAND2_2043(II10927,II10929,II10930);
  nand NAND2_2044(II10935,WX3355,II10927);
  nand NAND2_2045(II10936,WX3355,II10935);
  nand NAND2_2046(II10937,II10927,II10935);
  nand NAND2_2047(II10926,II10936,II10937);
  nand NAND2_2048(II10943,WX3419,WX3483);
  nand NAND2_2049(II10944,WX3419,II10943);
  nand NAND2_2050(II10945,WX3483,II10943);
  nand NAND2_2051(II10942,II10944,II10945);
  nand NAND2_2052(II10950,II10926,II10942);
  nand NAND2_2053(II10951,II10926,II10950);
  nand NAND2_2054(II10952,II10942,II10950);
  nand NAND2_2055(WX3516,II10951,II10952);
  nand NAND2_2056(II10959,WX3588,WX3293);
  nand NAND2_2057(II10960,WX3588,II10959);
  nand NAND2_2058(II10961,WX3293,II10959);
  nand NAND2_2059(II10958,II10960,II10961);
  nand NAND2_2060(II10966,WX3357,II10958);
  nand NAND2_2061(II10967,WX3357,II10966);
  nand NAND2_2062(II10968,II10958,II10966);
  nand NAND2_2063(II10957,II10967,II10968);
  nand NAND2_2064(II10974,WX3421,WX3485);
  nand NAND2_2065(II10975,WX3421,II10974);
  nand NAND2_2066(II10976,WX3485,II10974);
  nand NAND2_2067(II10973,II10975,II10976);
  nand NAND2_2068(II10981,II10957,II10973);
  nand NAND2_2069(II10982,II10957,II10981);
  nand NAND2_2070(II10983,II10973,II10981);
  nand NAND2_2071(WX3517,II10982,II10983);
  nand NAND2_2072(II11062,WX3166,WX3071);
  nand NAND2_2073(II11063,WX3166,II11062);
  nand NAND2_2074(II11064,WX3071,II11062);
  nand NAND2_2075(WX3592,II11063,II11064);
  nand NAND2_2076(II11075,WX3167,WX3073);
  nand NAND2_2077(II11076,WX3167,II11075);
  nand NAND2_2078(II11077,WX3073,II11075);
  nand NAND2_2079(WX3599,II11076,II11077);
  nand NAND2_2080(II11088,WX3168,WX3075);
  nand NAND2_2081(II11089,WX3168,II11088);
  nand NAND2_2082(II11090,WX3075,II11088);
  nand NAND2_2083(WX3606,II11089,II11090);
  nand NAND2_2084(II11101,WX3169,WX3077);
  nand NAND2_2085(II11102,WX3169,II11101);
  nand NAND2_2086(II11103,WX3077,II11101);
  nand NAND2_2087(WX3613,II11102,II11103);
  nand NAND2_2088(II11114,WX3170,WX3079);
  nand NAND2_2089(II11115,WX3170,II11114);
  nand NAND2_2090(II11116,WX3079,II11114);
  nand NAND2_2091(WX3620,II11115,II11116);
  nand NAND2_2092(II11127,WX3171,WX3081);
  nand NAND2_2093(II11128,WX3171,II11127);
  nand NAND2_2094(II11129,WX3081,II11127);
  nand NAND2_2095(WX3627,II11128,II11129);
  nand NAND2_2096(II11140,WX3172,WX3083);
  nand NAND2_2097(II11141,WX3172,II11140);
  nand NAND2_2098(II11142,WX3083,II11140);
  nand NAND2_2099(WX3634,II11141,II11142);
  nand NAND2_2100(II11153,WX3173,WX3085);
  nand NAND2_2101(II11154,WX3173,II11153);
  nand NAND2_2102(II11155,WX3085,II11153);
  nand NAND2_2103(WX3641,II11154,II11155);
  nand NAND2_2104(II11166,WX3174,WX3087);
  nand NAND2_2105(II11167,WX3174,II11166);
  nand NAND2_2106(II11168,WX3087,II11166);
  nand NAND2_2107(WX3648,II11167,II11168);
  nand NAND2_2108(II11179,WX3175,WX3089);
  nand NAND2_2109(II11180,WX3175,II11179);
  nand NAND2_2110(II11181,WX3089,II11179);
  nand NAND2_2111(WX3655,II11180,II11181);
  nand NAND2_2112(II11192,WX3176,WX3091);
  nand NAND2_2113(II11193,WX3176,II11192);
  nand NAND2_2114(II11194,WX3091,II11192);
  nand NAND2_2115(WX3662,II11193,II11194);
  nand NAND2_2116(II11205,WX3177,WX3093);
  nand NAND2_2117(II11206,WX3177,II11205);
  nand NAND2_2118(II11207,WX3093,II11205);
  nand NAND2_2119(WX3669,II11206,II11207);
  nand NAND2_2120(II11218,WX3178,WX3095);
  nand NAND2_2121(II11219,WX3178,II11218);
  nand NAND2_2122(II11220,WX3095,II11218);
  nand NAND2_2123(WX3676,II11219,II11220);
  nand NAND2_2124(II11231,WX3179,WX3097);
  nand NAND2_2125(II11232,WX3179,II11231);
  nand NAND2_2126(II11233,WX3097,II11231);
  nand NAND2_2127(WX3683,II11232,II11233);
  nand NAND2_2128(II11244,WX3180,WX3099);
  nand NAND2_2129(II11245,WX3180,II11244);
  nand NAND2_2130(II11246,WX3099,II11244);
  nand NAND2_2131(WX3690,II11245,II11246);
  nand NAND2_2132(II11257,WX3181,WX3101);
  nand NAND2_2133(II11258,WX3181,II11257);
  nand NAND2_2134(II11259,WX3101,II11257);
  nand NAND2_2135(WX3697,II11258,II11259);
  nand NAND2_2136(II11270,WX3182,WX3103);
  nand NAND2_2137(II11271,WX3182,II11270);
  nand NAND2_2138(II11272,WX3103,II11270);
  nand NAND2_2139(WX3704,II11271,II11272);
  nand NAND2_2140(II11283,WX3183,WX3105);
  nand NAND2_2141(II11284,WX3183,II11283);
  nand NAND2_2142(II11285,WX3105,II11283);
  nand NAND2_2143(WX3711,II11284,II11285);
  nand NAND2_2144(II11296,WX3184,WX3107);
  nand NAND2_2145(II11297,WX3184,II11296);
  nand NAND2_2146(II11298,WX3107,II11296);
  nand NAND2_2147(WX3718,II11297,II11298);
  nand NAND2_2148(II11309,WX3185,WX3109);
  nand NAND2_2149(II11310,WX3185,II11309);
  nand NAND2_2150(II11311,WX3109,II11309);
  nand NAND2_2151(WX3725,II11310,II11311);
  nand NAND2_2152(II11322,WX3186,WX3111);
  nand NAND2_2153(II11323,WX3186,II11322);
  nand NAND2_2154(II11324,WX3111,II11322);
  nand NAND2_2155(WX3732,II11323,II11324);
  nand NAND2_2156(II11335,WX3187,WX3113);
  nand NAND2_2157(II11336,WX3187,II11335);
  nand NAND2_2158(II11337,WX3113,II11335);
  nand NAND2_2159(WX3739,II11336,II11337);
  nand NAND2_2160(II11348,WX3188,WX3115);
  nand NAND2_2161(II11349,WX3188,II11348);
  nand NAND2_2162(II11350,WX3115,II11348);
  nand NAND2_2163(WX3746,II11349,II11350);
  nand NAND2_2164(II11361,WX3189,WX3117);
  nand NAND2_2165(II11362,WX3189,II11361);
  nand NAND2_2166(II11363,WX3117,II11361);
  nand NAND2_2167(WX3753,II11362,II11363);
  nand NAND2_2168(II11374,WX3190,WX3119);
  nand NAND2_2169(II11375,WX3190,II11374);
  nand NAND2_2170(II11376,WX3119,II11374);
  nand NAND2_2171(WX3760,II11375,II11376);
  nand NAND2_2172(II11387,WX3191,WX3121);
  nand NAND2_2173(II11388,WX3191,II11387);
  nand NAND2_2174(II11389,WX3121,II11387);
  nand NAND2_2175(WX3767,II11388,II11389);
  nand NAND2_2176(II11400,WX3192,WX3123);
  nand NAND2_2177(II11401,WX3192,II11400);
  nand NAND2_2178(II11402,WX3123,II11400);
  nand NAND2_2179(WX3774,II11401,II11402);
  nand NAND2_2180(II11413,WX3193,WX3125);
  nand NAND2_2181(II11414,WX3193,II11413);
  nand NAND2_2182(II11415,WX3125,II11413);
  nand NAND2_2183(WX3781,II11414,II11415);
  nand NAND2_2184(II11426,WX3194,WX3127);
  nand NAND2_2185(II11427,WX3194,II11426);
  nand NAND2_2186(II11428,WX3127,II11426);
  nand NAND2_2187(WX3788,II11427,II11428);
  nand NAND2_2188(II11439,WX3195,WX3129);
  nand NAND2_2189(II11440,WX3195,II11439);
  nand NAND2_2190(II11441,WX3129,II11439);
  nand NAND2_2191(WX3795,II11440,II11441);
  nand NAND2_2192(II11452,WX3196,WX3131);
  nand NAND2_2193(II11453,WX3196,II11452);
  nand NAND2_2194(II11454,WX3131,II11452);
  nand NAND2_2195(WX3802,II11453,II11454);
  nand NAND2_2196(II11465,WX3197,WX3133);
  nand NAND2_2197(II11466,WX3197,II11465);
  nand NAND2_2198(II11467,WX3133,II11465);
  nand NAND2_2199(WX3809,II11466,II11467);
  nand NAND2_2200(II11480,WX3213,CRC_OUT_7_31);
  nand NAND2_2201(II11481,WX3213,II11480);
  nand NAND2_2202(II11482,CRC_OUT_7_31,II11480);
  nand NAND2_2203(II11479,II11481,II11482);
  nand NAND2_2204(II11487,CRC_OUT_7_15,II11479);
  nand NAND2_2205(II11488,CRC_OUT_7_15,II11487);
  nand NAND2_2206(II11489,II11479,II11487);
  nand NAND2_2207(WX3817,II11488,II11489);
  nand NAND2_2208(II11495,WX3218,CRC_OUT_7_31);
  nand NAND2_2209(II11496,WX3218,II11495);
  nand NAND2_2210(II11497,CRC_OUT_7_31,II11495);
  nand NAND2_2211(II11494,II11496,II11497);
  nand NAND2_2212(II11502,CRC_OUT_7_10,II11494);
  nand NAND2_2213(II11503,CRC_OUT_7_10,II11502);
  nand NAND2_2214(II11504,II11494,II11502);
  nand NAND2_2215(WX3818,II11503,II11504);
  nand NAND2_2216(II11510,WX3225,CRC_OUT_7_31);
  nand NAND2_2217(II11511,WX3225,II11510);
  nand NAND2_2218(II11512,CRC_OUT_7_31,II11510);
  nand NAND2_2219(II11509,II11511,II11512);
  nand NAND2_2220(II11517,CRC_OUT_7_3,II11509);
  nand NAND2_2221(II11518,CRC_OUT_7_3,II11517);
  nand NAND2_2222(II11519,II11509,II11517);
  nand NAND2_2223(WX3819,II11518,II11519);
  nand NAND2_2224(II11524,WX3229,CRC_OUT_7_31);
  nand NAND2_2225(II11525,WX3229,II11524);
  nand NAND2_2226(II11526,CRC_OUT_7_31,II11524);
  nand NAND2_2227(WX3820,II11525,II11526);
  nand NAND2_2228(II11531,WX3198,CRC_OUT_7_30);
  nand NAND2_2229(II11532,WX3198,II11531);
  nand NAND2_2230(II11533,CRC_OUT_7_30,II11531);
  nand NAND2_2231(WX3821,II11532,II11533);
  nand NAND2_2232(II11538,WX3199,CRC_OUT_7_29);
  nand NAND2_2233(II11539,WX3199,II11538);
  nand NAND2_2234(II11540,CRC_OUT_7_29,II11538);
  nand NAND2_2235(WX3822,II11539,II11540);
  nand NAND2_2236(II11545,WX3200,CRC_OUT_7_28);
  nand NAND2_2237(II11546,WX3200,II11545);
  nand NAND2_2238(II11547,CRC_OUT_7_28,II11545);
  nand NAND2_2239(WX3823,II11546,II11547);
  nand NAND2_2240(II11552,WX3201,CRC_OUT_7_27);
  nand NAND2_2241(II11553,WX3201,II11552);
  nand NAND2_2242(II11554,CRC_OUT_7_27,II11552);
  nand NAND2_2243(WX3824,II11553,II11554);
  nand NAND2_2244(II11559,WX3202,CRC_OUT_7_26);
  nand NAND2_2245(II11560,WX3202,II11559);
  nand NAND2_2246(II11561,CRC_OUT_7_26,II11559);
  nand NAND2_2247(WX3825,II11560,II11561);
  nand NAND2_2248(II11566,WX3203,CRC_OUT_7_25);
  nand NAND2_2249(II11567,WX3203,II11566);
  nand NAND2_2250(II11568,CRC_OUT_7_25,II11566);
  nand NAND2_2251(WX3826,II11567,II11568);
  nand NAND2_2252(II11573,WX3204,CRC_OUT_7_24);
  nand NAND2_2253(II11574,WX3204,II11573);
  nand NAND2_2254(II11575,CRC_OUT_7_24,II11573);
  nand NAND2_2255(WX3827,II11574,II11575);
  nand NAND2_2256(II11580,WX3205,CRC_OUT_7_23);
  nand NAND2_2257(II11581,WX3205,II11580);
  nand NAND2_2258(II11582,CRC_OUT_7_23,II11580);
  nand NAND2_2259(WX3828,II11581,II11582);
  nand NAND2_2260(II11587,WX3206,CRC_OUT_7_22);
  nand NAND2_2261(II11588,WX3206,II11587);
  nand NAND2_2262(II11589,CRC_OUT_7_22,II11587);
  nand NAND2_2263(WX3829,II11588,II11589);
  nand NAND2_2264(II11594,WX3207,CRC_OUT_7_21);
  nand NAND2_2265(II11595,WX3207,II11594);
  nand NAND2_2266(II11596,CRC_OUT_7_21,II11594);
  nand NAND2_2267(WX3830,II11595,II11596);
  nand NAND2_2268(II11601,WX3208,CRC_OUT_7_20);
  nand NAND2_2269(II11602,WX3208,II11601);
  nand NAND2_2270(II11603,CRC_OUT_7_20,II11601);
  nand NAND2_2271(WX3831,II11602,II11603);
  nand NAND2_2272(II11608,WX3209,CRC_OUT_7_19);
  nand NAND2_2273(II11609,WX3209,II11608);
  nand NAND2_2274(II11610,CRC_OUT_7_19,II11608);
  nand NAND2_2275(WX3832,II11609,II11610);
  nand NAND2_2276(II11615,WX3210,CRC_OUT_7_18);
  nand NAND2_2277(II11616,WX3210,II11615);
  nand NAND2_2278(II11617,CRC_OUT_7_18,II11615);
  nand NAND2_2279(WX3833,II11616,II11617);
  nand NAND2_2280(II11622,WX3211,CRC_OUT_7_17);
  nand NAND2_2281(II11623,WX3211,II11622);
  nand NAND2_2282(II11624,CRC_OUT_7_17,II11622);
  nand NAND2_2283(WX3834,II11623,II11624);
  nand NAND2_2284(II11629,WX3212,CRC_OUT_7_16);
  nand NAND2_2285(II11630,WX3212,II11629);
  nand NAND2_2286(II11631,CRC_OUT_7_16,II11629);
  nand NAND2_2287(WX3835,II11630,II11631);
  nand NAND2_2288(II11636,WX3214,CRC_OUT_7_14);
  nand NAND2_2289(II11637,WX3214,II11636);
  nand NAND2_2290(II11638,CRC_OUT_7_14,II11636);
  nand NAND2_2291(WX3836,II11637,II11638);
  nand NAND2_2292(II11643,WX3215,CRC_OUT_7_13);
  nand NAND2_2293(II11644,WX3215,II11643);
  nand NAND2_2294(II11645,CRC_OUT_7_13,II11643);
  nand NAND2_2295(WX3837,II11644,II11645);
  nand NAND2_2296(II11650,WX3216,CRC_OUT_7_12);
  nand NAND2_2297(II11651,WX3216,II11650);
  nand NAND2_2298(II11652,CRC_OUT_7_12,II11650);
  nand NAND2_2299(WX3838,II11651,II11652);
  nand NAND2_2300(II11657,WX3217,CRC_OUT_7_11);
  nand NAND2_2301(II11658,WX3217,II11657);
  nand NAND2_2302(II11659,CRC_OUT_7_11,II11657);
  nand NAND2_2303(WX3839,II11658,II11659);
  nand NAND2_2304(II11664,WX3219,CRC_OUT_7_9);
  nand NAND2_2305(II11665,WX3219,II11664);
  nand NAND2_2306(II11666,CRC_OUT_7_9,II11664);
  nand NAND2_2307(WX3840,II11665,II11666);
  nand NAND2_2308(II11671,WX3220,CRC_OUT_7_8);
  nand NAND2_2309(II11672,WX3220,II11671);
  nand NAND2_2310(II11673,CRC_OUT_7_8,II11671);
  nand NAND2_2311(WX3841,II11672,II11673);
  nand NAND2_2312(II11678,WX3221,CRC_OUT_7_7);
  nand NAND2_2313(II11679,WX3221,II11678);
  nand NAND2_2314(II11680,CRC_OUT_7_7,II11678);
  nand NAND2_2315(WX3842,II11679,II11680);
  nand NAND2_2316(II11685,WX3222,CRC_OUT_7_6);
  nand NAND2_2317(II11686,WX3222,II11685);
  nand NAND2_2318(II11687,CRC_OUT_7_6,II11685);
  nand NAND2_2319(WX3843,II11686,II11687);
  nand NAND2_2320(II11692,WX3223,CRC_OUT_7_5);
  nand NAND2_2321(II11693,WX3223,II11692);
  nand NAND2_2322(II11694,CRC_OUT_7_5,II11692);
  nand NAND2_2323(WX3844,II11693,II11694);
  nand NAND2_2324(II11699,WX3224,CRC_OUT_7_4);
  nand NAND2_2325(II11700,WX3224,II11699);
  nand NAND2_2326(II11701,CRC_OUT_7_4,II11699);
  nand NAND2_2327(WX3845,II11700,II11701);
  nand NAND2_2328(II11706,WX3226,CRC_OUT_7_2);
  nand NAND2_2329(II11707,WX3226,II11706);
  nand NAND2_2330(II11708,CRC_OUT_7_2,II11706);
  nand NAND2_2331(WX3846,II11707,II11708);
  nand NAND2_2332(II11713,WX3227,CRC_OUT_7_1);
  nand NAND2_2333(II11714,WX3227,II11713);
  nand NAND2_2334(II11715,CRC_OUT_7_1,II11713);
  nand NAND2_2335(WX3847,II11714,II11715);
  nand NAND2_2336(II11720,WX3228,CRC_OUT_7_0);
  nand NAND2_2337(II11721,WX3228,II11720);
  nand NAND2_2338(II11722,CRC_OUT_7_0,II11720);
  nand NAND2_2339(WX3848,II11721,II11722);
  nand NAND2_2340(II14003,WX4880,WX4524);
  nand NAND2_2341(II14004,WX4880,II14003);
  nand NAND2_2342(II14005,WX4524,II14003);
  nand NAND2_2343(II14002,II14004,II14005);
  nand NAND2_2344(II14010,WX4588,II14002);
  nand NAND2_2345(II14011,WX4588,II14010);
  nand NAND2_2346(II14012,II14002,II14010);
  nand NAND2_2347(II14001,II14011,II14012);
  nand NAND2_2348(II14018,WX4652,WX4716);
  nand NAND2_2349(II14019,WX4652,II14018);
  nand NAND2_2350(II14020,WX4716,II14018);
  nand NAND2_2351(II14017,II14019,II14020);
  nand NAND2_2352(II14025,II14001,II14017);
  nand NAND2_2353(II14026,II14001,II14025);
  nand NAND2_2354(II14027,II14017,II14025);
  nand NAND2_2355(WX4779,II14026,II14027);
  nand NAND2_2356(II14034,WX4880,WX4526);
  nand NAND2_2357(II14035,WX4880,II14034);
  nand NAND2_2358(II14036,WX4526,II14034);
  nand NAND2_2359(II14033,II14035,II14036);
  nand NAND2_2360(II14041,WX4590,II14033);
  nand NAND2_2361(II14042,WX4590,II14041);
  nand NAND2_2362(II14043,II14033,II14041);
  nand NAND2_2363(II14032,II14042,II14043);
  nand NAND2_2364(II14049,WX4654,WX4718);
  nand NAND2_2365(II14050,WX4654,II14049);
  nand NAND2_2366(II14051,WX4718,II14049);
  nand NAND2_2367(II14048,II14050,II14051);
  nand NAND2_2368(II14056,II14032,II14048);
  nand NAND2_2369(II14057,II14032,II14056);
  nand NAND2_2370(II14058,II14048,II14056);
  nand NAND2_2371(WX4780,II14057,II14058);
  nand NAND2_2372(II14065,WX4880,WX4528);
  nand NAND2_2373(II14066,WX4880,II14065);
  nand NAND2_2374(II14067,WX4528,II14065);
  nand NAND2_2375(II14064,II14066,II14067);
  nand NAND2_2376(II14072,WX4592,II14064);
  nand NAND2_2377(II14073,WX4592,II14072);
  nand NAND2_2378(II14074,II14064,II14072);
  nand NAND2_2379(II14063,II14073,II14074);
  nand NAND2_2380(II14080,WX4656,WX4720);
  nand NAND2_2381(II14081,WX4656,II14080);
  nand NAND2_2382(II14082,WX4720,II14080);
  nand NAND2_2383(II14079,II14081,II14082);
  nand NAND2_2384(II14087,II14063,II14079);
  nand NAND2_2385(II14088,II14063,II14087);
  nand NAND2_2386(II14089,II14079,II14087);
  nand NAND2_2387(WX4781,II14088,II14089);
  nand NAND2_2388(II14096,WX4880,WX4530);
  nand NAND2_2389(II14097,WX4880,II14096);
  nand NAND2_2390(II14098,WX4530,II14096);
  nand NAND2_2391(II14095,II14097,II14098);
  nand NAND2_2392(II14103,WX4594,II14095);
  nand NAND2_2393(II14104,WX4594,II14103);
  nand NAND2_2394(II14105,II14095,II14103);
  nand NAND2_2395(II14094,II14104,II14105);
  nand NAND2_2396(II14111,WX4658,WX4722);
  nand NAND2_2397(II14112,WX4658,II14111);
  nand NAND2_2398(II14113,WX4722,II14111);
  nand NAND2_2399(II14110,II14112,II14113);
  nand NAND2_2400(II14118,II14094,II14110);
  nand NAND2_2401(II14119,II14094,II14118);
  nand NAND2_2402(II14120,II14110,II14118);
  nand NAND2_2403(WX4782,II14119,II14120);
  nand NAND2_2404(II14127,WX4880,WX4532);
  nand NAND2_2405(II14128,WX4880,II14127);
  nand NAND2_2406(II14129,WX4532,II14127);
  nand NAND2_2407(II14126,II14128,II14129);
  nand NAND2_2408(II14134,WX4596,II14126);
  nand NAND2_2409(II14135,WX4596,II14134);
  nand NAND2_2410(II14136,II14126,II14134);
  nand NAND2_2411(II14125,II14135,II14136);
  nand NAND2_2412(II14142,WX4660,WX4724);
  nand NAND2_2413(II14143,WX4660,II14142);
  nand NAND2_2414(II14144,WX4724,II14142);
  nand NAND2_2415(II14141,II14143,II14144);
  nand NAND2_2416(II14149,II14125,II14141);
  nand NAND2_2417(II14150,II14125,II14149);
  nand NAND2_2418(II14151,II14141,II14149);
  nand NAND2_2419(WX4783,II14150,II14151);
  nand NAND2_2420(II14158,WX4880,WX4534);
  nand NAND2_2421(II14159,WX4880,II14158);
  nand NAND2_2422(II14160,WX4534,II14158);
  nand NAND2_2423(II14157,II14159,II14160);
  nand NAND2_2424(II14165,WX4598,II14157);
  nand NAND2_2425(II14166,WX4598,II14165);
  nand NAND2_2426(II14167,II14157,II14165);
  nand NAND2_2427(II14156,II14166,II14167);
  nand NAND2_2428(II14173,WX4662,WX4726);
  nand NAND2_2429(II14174,WX4662,II14173);
  nand NAND2_2430(II14175,WX4726,II14173);
  nand NAND2_2431(II14172,II14174,II14175);
  nand NAND2_2432(II14180,II14156,II14172);
  nand NAND2_2433(II14181,II14156,II14180);
  nand NAND2_2434(II14182,II14172,II14180);
  nand NAND2_2435(WX4784,II14181,II14182);
  nand NAND2_2436(II14189,WX4880,WX4536);
  nand NAND2_2437(II14190,WX4880,II14189);
  nand NAND2_2438(II14191,WX4536,II14189);
  nand NAND2_2439(II14188,II14190,II14191);
  nand NAND2_2440(II14196,WX4600,II14188);
  nand NAND2_2441(II14197,WX4600,II14196);
  nand NAND2_2442(II14198,II14188,II14196);
  nand NAND2_2443(II14187,II14197,II14198);
  nand NAND2_2444(II14204,WX4664,WX4728);
  nand NAND2_2445(II14205,WX4664,II14204);
  nand NAND2_2446(II14206,WX4728,II14204);
  nand NAND2_2447(II14203,II14205,II14206);
  nand NAND2_2448(II14211,II14187,II14203);
  nand NAND2_2449(II14212,II14187,II14211);
  nand NAND2_2450(II14213,II14203,II14211);
  nand NAND2_2451(WX4785,II14212,II14213);
  nand NAND2_2452(II14220,WX4880,WX4538);
  nand NAND2_2453(II14221,WX4880,II14220);
  nand NAND2_2454(II14222,WX4538,II14220);
  nand NAND2_2455(II14219,II14221,II14222);
  nand NAND2_2456(II14227,WX4602,II14219);
  nand NAND2_2457(II14228,WX4602,II14227);
  nand NAND2_2458(II14229,II14219,II14227);
  nand NAND2_2459(II14218,II14228,II14229);
  nand NAND2_2460(II14235,WX4666,WX4730);
  nand NAND2_2461(II14236,WX4666,II14235);
  nand NAND2_2462(II14237,WX4730,II14235);
  nand NAND2_2463(II14234,II14236,II14237);
  nand NAND2_2464(II14242,II14218,II14234);
  nand NAND2_2465(II14243,II14218,II14242);
  nand NAND2_2466(II14244,II14234,II14242);
  nand NAND2_2467(WX4786,II14243,II14244);
  nand NAND2_2468(II14251,WX4880,WX4540);
  nand NAND2_2469(II14252,WX4880,II14251);
  nand NAND2_2470(II14253,WX4540,II14251);
  nand NAND2_2471(II14250,II14252,II14253);
  nand NAND2_2472(II14258,WX4604,II14250);
  nand NAND2_2473(II14259,WX4604,II14258);
  nand NAND2_2474(II14260,II14250,II14258);
  nand NAND2_2475(II14249,II14259,II14260);
  nand NAND2_2476(II14266,WX4668,WX4732);
  nand NAND2_2477(II14267,WX4668,II14266);
  nand NAND2_2478(II14268,WX4732,II14266);
  nand NAND2_2479(II14265,II14267,II14268);
  nand NAND2_2480(II14273,II14249,II14265);
  nand NAND2_2481(II14274,II14249,II14273);
  nand NAND2_2482(II14275,II14265,II14273);
  nand NAND2_2483(WX4787,II14274,II14275);
  nand NAND2_2484(II14282,WX4880,WX4542);
  nand NAND2_2485(II14283,WX4880,II14282);
  nand NAND2_2486(II14284,WX4542,II14282);
  nand NAND2_2487(II14281,II14283,II14284);
  nand NAND2_2488(II14289,WX4606,II14281);
  nand NAND2_2489(II14290,WX4606,II14289);
  nand NAND2_2490(II14291,II14281,II14289);
  nand NAND2_2491(II14280,II14290,II14291);
  nand NAND2_2492(II14297,WX4670,WX4734);
  nand NAND2_2493(II14298,WX4670,II14297);
  nand NAND2_2494(II14299,WX4734,II14297);
  nand NAND2_2495(II14296,II14298,II14299);
  nand NAND2_2496(II14304,II14280,II14296);
  nand NAND2_2497(II14305,II14280,II14304);
  nand NAND2_2498(II14306,II14296,II14304);
  nand NAND2_2499(WX4788,II14305,II14306);
  nand NAND2_2500(II14313,WX4880,WX4544);
  nand NAND2_2501(II14314,WX4880,II14313);
  nand NAND2_2502(II14315,WX4544,II14313);
  nand NAND2_2503(II14312,II14314,II14315);
  nand NAND2_2504(II14320,WX4608,II14312);
  nand NAND2_2505(II14321,WX4608,II14320);
  nand NAND2_2506(II14322,II14312,II14320);
  nand NAND2_2507(II14311,II14321,II14322);
  nand NAND2_2508(II14328,WX4672,WX4736);
  nand NAND2_2509(II14329,WX4672,II14328);
  nand NAND2_2510(II14330,WX4736,II14328);
  nand NAND2_2511(II14327,II14329,II14330);
  nand NAND2_2512(II14335,II14311,II14327);
  nand NAND2_2513(II14336,II14311,II14335);
  nand NAND2_2514(II14337,II14327,II14335);
  nand NAND2_2515(WX4789,II14336,II14337);
  nand NAND2_2516(II14344,WX4880,WX4546);
  nand NAND2_2517(II14345,WX4880,II14344);
  nand NAND2_2518(II14346,WX4546,II14344);
  nand NAND2_2519(II14343,II14345,II14346);
  nand NAND2_2520(II14351,WX4610,II14343);
  nand NAND2_2521(II14352,WX4610,II14351);
  nand NAND2_2522(II14353,II14343,II14351);
  nand NAND2_2523(II14342,II14352,II14353);
  nand NAND2_2524(II14359,WX4674,WX4738);
  nand NAND2_2525(II14360,WX4674,II14359);
  nand NAND2_2526(II14361,WX4738,II14359);
  nand NAND2_2527(II14358,II14360,II14361);
  nand NAND2_2528(II14366,II14342,II14358);
  nand NAND2_2529(II14367,II14342,II14366);
  nand NAND2_2530(II14368,II14358,II14366);
  nand NAND2_2531(WX4790,II14367,II14368);
  nand NAND2_2532(II14375,WX4880,WX4548);
  nand NAND2_2533(II14376,WX4880,II14375);
  nand NAND2_2534(II14377,WX4548,II14375);
  nand NAND2_2535(II14374,II14376,II14377);
  nand NAND2_2536(II14382,WX4612,II14374);
  nand NAND2_2537(II14383,WX4612,II14382);
  nand NAND2_2538(II14384,II14374,II14382);
  nand NAND2_2539(II14373,II14383,II14384);
  nand NAND2_2540(II14390,WX4676,WX4740);
  nand NAND2_2541(II14391,WX4676,II14390);
  nand NAND2_2542(II14392,WX4740,II14390);
  nand NAND2_2543(II14389,II14391,II14392);
  nand NAND2_2544(II14397,II14373,II14389);
  nand NAND2_2545(II14398,II14373,II14397);
  nand NAND2_2546(II14399,II14389,II14397);
  nand NAND2_2547(WX4791,II14398,II14399);
  nand NAND2_2548(II14406,WX4880,WX4550);
  nand NAND2_2549(II14407,WX4880,II14406);
  nand NAND2_2550(II14408,WX4550,II14406);
  nand NAND2_2551(II14405,II14407,II14408);
  nand NAND2_2552(II14413,WX4614,II14405);
  nand NAND2_2553(II14414,WX4614,II14413);
  nand NAND2_2554(II14415,II14405,II14413);
  nand NAND2_2555(II14404,II14414,II14415);
  nand NAND2_2556(II14421,WX4678,WX4742);
  nand NAND2_2557(II14422,WX4678,II14421);
  nand NAND2_2558(II14423,WX4742,II14421);
  nand NAND2_2559(II14420,II14422,II14423);
  nand NAND2_2560(II14428,II14404,II14420);
  nand NAND2_2561(II14429,II14404,II14428);
  nand NAND2_2562(II14430,II14420,II14428);
  nand NAND2_2563(WX4792,II14429,II14430);
  nand NAND2_2564(II14437,WX4880,WX4552);
  nand NAND2_2565(II14438,WX4880,II14437);
  nand NAND2_2566(II14439,WX4552,II14437);
  nand NAND2_2567(II14436,II14438,II14439);
  nand NAND2_2568(II14444,WX4616,II14436);
  nand NAND2_2569(II14445,WX4616,II14444);
  nand NAND2_2570(II14446,II14436,II14444);
  nand NAND2_2571(II14435,II14445,II14446);
  nand NAND2_2572(II14452,WX4680,WX4744);
  nand NAND2_2573(II14453,WX4680,II14452);
  nand NAND2_2574(II14454,WX4744,II14452);
  nand NAND2_2575(II14451,II14453,II14454);
  nand NAND2_2576(II14459,II14435,II14451);
  nand NAND2_2577(II14460,II14435,II14459);
  nand NAND2_2578(II14461,II14451,II14459);
  nand NAND2_2579(WX4793,II14460,II14461);
  nand NAND2_2580(II14468,WX4880,WX4554);
  nand NAND2_2581(II14469,WX4880,II14468);
  nand NAND2_2582(II14470,WX4554,II14468);
  nand NAND2_2583(II14467,II14469,II14470);
  nand NAND2_2584(II14475,WX4618,II14467);
  nand NAND2_2585(II14476,WX4618,II14475);
  nand NAND2_2586(II14477,II14467,II14475);
  nand NAND2_2587(II14466,II14476,II14477);
  nand NAND2_2588(II14483,WX4682,WX4746);
  nand NAND2_2589(II14484,WX4682,II14483);
  nand NAND2_2590(II14485,WX4746,II14483);
  nand NAND2_2591(II14482,II14484,II14485);
  nand NAND2_2592(II14490,II14466,II14482);
  nand NAND2_2593(II14491,II14466,II14490);
  nand NAND2_2594(II14492,II14482,II14490);
  nand NAND2_2595(WX4794,II14491,II14492);
  nand NAND2_2596(II14499,WX4881,WX4556);
  nand NAND2_2597(II14500,WX4881,II14499);
  nand NAND2_2598(II14501,WX4556,II14499);
  nand NAND2_2599(II14498,II14500,II14501);
  nand NAND2_2600(II14506,WX4620,II14498);
  nand NAND2_2601(II14507,WX4620,II14506);
  nand NAND2_2602(II14508,II14498,II14506);
  nand NAND2_2603(II14497,II14507,II14508);
  nand NAND2_2604(II14514,WX4684,WX4748);
  nand NAND2_2605(II14515,WX4684,II14514);
  nand NAND2_2606(II14516,WX4748,II14514);
  nand NAND2_2607(II14513,II14515,II14516);
  nand NAND2_2608(II14521,II14497,II14513);
  nand NAND2_2609(II14522,II14497,II14521);
  nand NAND2_2610(II14523,II14513,II14521);
  nand NAND2_2611(WX4795,II14522,II14523);
  nand NAND2_2612(II14530,WX4881,WX4558);
  nand NAND2_2613(II14531,WX4881,II14530);
  nand NAND2_2614(II14532,WX4558,II14530);
  nand NAND2_2615(II14529,II14531,II14532);
  nand NAND2_2616(II14537,WX4622,II14529);
  nand NAND2_2617(II14538,WX4622,II14537);
  nand NAND2_2618(II14539,II14529,II14537);
  nand NAND2_2619(II14528,II14538,II14539);
  nand NAND2_2620(II14545,WX4686,WX4750);
  nand NAND2_2621(II14546,WX4686,II14545);
  nand NAND2_2622(II14547,WX4750,II14545);
  nand NAND2_2623(II14544,II14546,II14547);
  nand NAND2_2624(II14552,II14528,II14544);
  nand NAND2_2625(II14553,II14528,II14552);
  nand NAND2_2626(II14554,II14544,II14552);
  nand NAND2_2627(WX4796,II14553,II14554);
  nand NAND2_2628(II14561,WX4881,WX4560);
  nand NAND2_2629(II14562,WX4881,II14561);
  nand NAND2_2630(II14563,WX4560,II14561);
  nand NAND2_2631(II14560,II14562,II14563);
  nand NAND2_2632(II14568,WX4624,II14560);
  nand NAND2_2633(II14569,WX4624,II14568);
  nand NAND2_2634(II14570,II14560,II14568);
  nand NAND2_2635(II14559,II14569,II14570);
  nand NAND2_2636(II14576,WX4688,WX4752);
  nand NAND2_2637(II14577,WX4688,II14576);
  nand NAND2_2638(II14578,WX4752,II14576);
  nand NAND2_2639(II14575,II14577,II14578);
  nand NAND2_2640(II14583,II14559,II14575);
  nand NAND2_2641(II14584,II14559,II14583);
  nand NAND2_2642(II14585,II14575,II14583);
  nand NAND2_2643(WX4797,II14584,II14585);
  nand NAND2_2644(II14592,WX4881,WX4562);
  nand NAND2_2645(II14593,WX4881,II14592);
  nand NAND2_2646(II14594,WX4562,II14592);
  nand NAND2_2647(II14591,II14593,II14594);
  nand NAND2_2648(II14599,WX4626,II14591);
  nand NAND2_2649(II14600,WX4626,II14599);
  nand NAND2_2650(II14601,II14591,II14599);
  nand NAND2_2651(II14590,II14600,II14601);
  nand NAND2_2652(II14607,WX4690,WX4754);
  nand NAND2_2653(II14608,WX4690,II14607);
  nand NAND2_2654(II14609,WX4754,II14607);
  nand NAND2_2655(II14606,II14608,II14609);
  nand NAND2_2656(II14614,II14590,II14606);
  nand NAND2_2657(II14615,II14590,II14614);
  nand NAND2_2658(II14616,II14606,II14614);
  nand NAND2_2659(WX4798,II14615,II14616);
  nand NAND2_2660(II14623,WX4881,WX4564);
  nand NAND2_2661(II14624,WX4881,II14623);
  nand NAND2_2662(II14625,WX4564,II14623);
  nand NAND2_2663(II14622,II14624,II14625);
  nand NAND2_2664(II14630,WX4628,II14622);
  nand NAND2_2665(II14631,WX4628,II14630);
  nand NAND2_2666(II14632,II14622,II14630);
  nand NAND2_2667(II14621,II14631,II14632);
  nand NAND2_2668(II14638,WX4692,WX4756);
  nand NAND2_2669(II14639,WX4692,II14638);
  nand NAND2_2670(II14640,WX4756,II14638);
  nand NAND2_2671(II14637,II14639,II14640);
  nand NAND2_2672(II14645,II14621,II14637);
  nand NAND2_2673(II14646,II14621,II14645);
  nand NAND2_2674(II14647,II14637,II14645);
  nand NAND2_2675(WX4799,II14646,II14647);
  nand NAND2_2676(II14654,WX4881,WX4566);
  nand NAND2_2677(II14655,WX4881,II14654);
  nand NAND2_2678(II14656,WX4566,II14654);
  nand NAND2_2679(II14653,II14655,II14656);
  nand NAND2_2680(II14661,WX4630,II14653);
  nand NAND2_2681(II14662,WX4630,II14661);
  nand NAND2_2682(II14663,II14653,II14661);
  nand NAND2_2683(II14652,II14662,II14663);
  nand NAND2_2684(II14669,WX4694,WX4758);
  nand NAND2_2685(II14670,WX4694,II14669);
  nand NAND2_2686(II14671,WX4758,II14669);
  nand NAND2_2687(II14668,II14670,II14671);
  nand NAND2_2688(II14676,II14652,II14668);
  nand NAND2_2689(II14677,II14652,II14676);
  nand NAND2_2690(II14678,II14668,II14676);
  nand NAND2_2691(WX4800,II14677,II14678);
  nand NAND2_2692(II14685,WX4881,WX4568);
  nand NAND2_2693(II14686,WX4881,II14685);
  nand NAND2_2694(II14687,WX4568,II14685);
  nand NAND2_2695(II14684,II14686,II14687);
  nand NAND2_2696(II14692,WX4632,II14684);
  nand NAND2_2697(II14693,WX4632,II14692);
  nand NAND2_2698(II14694,II14684,II14692);
  nand NAND2_2699(II14683,II14693,II14694);
  nand NAND2_2700(II14700,WX4696,WX4760);
  nand NAND2_2701(II14701,WX4696,II14700);
  nand NAND2_2702(II14702,WX4760,II14700);
  nand NAND2_2703(II14699,II14701,II14702);
  nand NAND2_2704(II14707,II14683,II14699);
  nand NAND2_2705(II14708,II14683,II14707);
  nand NAND2_2706(II14709,II14699,II14707);
  nand NAND2_2707(WX4801,II14708,II14709);
  nand NAND2_2708(II14716,WX4881,WX4570);
  nand NAND2_2709(II14717,WX4881,II14716);
  nand NAND2_2710(II14718,WX4570,II14716);
  nand NAND2_2711(II14715,II14717,II14718);
  nand NAND2_2712(II14723,WX4634,II14715);
  nand NAND2_2713(II14724,WX4634,II14723);
  nand NAND2_2714(II14725,II14715,II14723);
  nand NAND2_2715(II14714,II14724,II14725);
  nand NAND2_2716(II14731,WX4698,WX4762);
  nand NAND2_2717(II14732,WX4698,II14731);
  nand NAND2_2718(II14733,WX4762,II14731);
  nand NAND2_2719(II14730,II14732,II14733);
  nand NAND2_2720(II14738,II14714,II14730);
  nand NAND2_2721(II14739,II14714,II14738);
  nand NAND2_2722(II14740,II14730,II14738);
  nand NAND2_2723(WX4802,II14739,II14740);
  nand NAND2_2724(II14747,WX4881,WX4572);
  nand NAND2_2725(II14748,WX4881,II14747);
  nand NAND2_2726(II14749,WX4572,II14747);
  nand NAND2_2727(II14746,II14748,II14749);
  nand NAND2_2728(II14754,WX4636,II14746);
  nand NAND2_2729(II14755,WX4636,II14754);
  nand NAND2_2730(II14756,II14746,II14754);
  nand NAND2_2731(II14745,II14755,II14756);
  nand NAND2_2732(II14762,WX4700,WX4764);
  nand NAND2_2733(II14763,WX4700,II14762);
  nand NAND2_2734(II14764,WX4764,II14762);
  nand NAND2_2735(II14761,II14763,II14764);
  nand NAND2_2736(II14769,II14745,II14761);
  nand NAND2_2737(II14770,II14745,II14769);
  nand NAND2_2738(II14771,II14761,II14769);
  nand NAND2_2739(WX4803,II14770,II14771);
  nand NAND2_2740(II14778,WX4881,WX4574);
  nand NAND2_2741(II14779,WX4881,II14778);
  nand NAND2_2742(II14780,WX4574,II14778);
  nand NAND2_2743(II14777,II14779,II14780);
  nand NAND2_2744(II14785,WX4638,II14777);
  nand NAND2_2745(II14786,WX4638,II14785);
  nand NAND2_2746(II14787,II14777,II14785);
  nand NAND2_2747(II14776,II14786,II14787);
  nand NAND2_2748(II14793,WX4702,WX4766);
  nand NAND2_2749(II14794,WX4702,II14793);
  nand NAND2_2750(II14795,WX4766,II14793);
  nand NAND2_2751(II14792,II14794,II14795);
  nand NAND2_2752(II14800,II14776,II14792);
  nand NAND2_2753(II14801,II14776,II14800);
  nand NAND2_2754(II14802,II14792,II14800);
  nand NAND2_2755(WX4804,II14801,II14802);
  nand NAND2_2756(II14809,WX4881,WX4576);
  nand NAND2_2757(II14810,WX4881,II14809);
  nand NAND2_2758(II14811,WX4576,II14809);
  nand NAND2_2759(II14808,II14810,II14811);
  nand NAND2_2760(II14816,WX4640,II14808);
  nand NAND2_2761(II14817,WX4640,II14816);
  nand NAND2_2762(II14818,II14808,II14816);
  nand NAND2_2763(II14807,II14817,II14818);
  nand NAND2_2764(II14824,WX4704,WX4768);
  nand NAND2_2765(II14825,WX4704,II14824);
  nand NAND2_2766(II14826,WX4768,II14824);
  nand NAND2_2767(II14823,II14825,II14826);
  nand NAND2_2768(II14831,II14807,II14823);
  nand NAND2_2769(II14832,II14807,II14831);
  nand NAND2_2770(II14833,II14823,II14831);
  nand NAND2_2771(WX4805,II14832,II14833);
  nand NAND2_2772(II14840,WX4881,WX4578);
  nand NAND2_2773(II14841,WX4881,II14840);
  nand NAND2_2774(II14842,WX4578,II14840);
  nand NAND2_2775(II14839,II14841,II14842);
  nand NAND2_2776(II14847,WX4642,II14839);
  nand NAND2_2777(II14848,WX4642,II14847);
  nand NAND2_2778(II14849,II14839,II14847);
  nand NAND2_2779(II14838,II14848,II14849);
  nand NAND2_2780(II14855,WX4706,WX4770);
  nand NAND2_2781(II14856,WX4706,II14855);
  nand NAND2_2782(II14857,WX4770,II14855);
  nand NAND2_2783(II14854,II14856,II14857);
  nand NAND2_2784(II14862,II14838,II14854);
  nand NAND2_2785(II14863,II14838,II14862);
  nand NAND2_2786(II14864,II14854,II14862);
  nand NAND2_2787(WX4806,II14863,II14864);
  nand NAND2_2788(II14871,WX4881,WX4580);
  nand NAND2_2789(II14872,WX4881,II14871);
  nand NAND2_2790(II14873,WX4580,II14871);
  nand NAND2_2791(II14870,II14872,II14873);
  nand NAND2_2792(II14878,WX4644,II14870);
  nand NAND2_2793(II14879,WX4644,II14878);
  nand NAND2_2794(II14880,II14870,II14878);
  nand NAND2_2795(II14869,II14879,II14880);
  nand NAND2_2796(II14886,WX4708,WX4772);
  nand NAND2_2797(II14887,WX4708,II14886);
  nand NAND2_2798(II14888,WX4772,II14886);
  nand NAND2_2799(II14885,II14887,II14888);
  nand NAND2_2800(II14893,II14869,II14885);
  nand NAND2_2801(II14894,II14869,II14893);
  nand NAND2_2802(II14895,II14885,II14893);
  nand NAND2_2803(WX4807,II14894,II14895);
  nand NAND2_2804(II14902,WX4881,WX4582);
  nand NAND2_2805(II14903,WX4881,II14902);
  nand NAND2_2806(II14904,WX4582,II14902);
  nand NAND2_2807(II14901,II14903,II14904);
  nand NAND2_2808(II14909,WX4646,II14901);
  nand NAND2_2809(II14910,WX4646,II14909);
  nand NAND2_2810(II14911,II14901,II14909);
  nand NAND2_2811(II14900,II14910,II14911);
  nand NAND2_2812(II14917,WX4710,WX4774);
  nand NAND2_2813(II14918,WX4710,II14917);
  nand NAND2_2814(II14919,WX4774,II14917);
  nand NAND2_2815(II14916,II14918,II14919);
  nand NAND2_2816(II14924,II14900,II14916);
  nand NAND2_2817(II14925,II14900,II14924);
  nand NAND2_2818(II14926,II14916,II14924);
  nand NAND2_2819(WX4808,II14925,II14926);
  nand NAND2_2820(II14933,WX4881,WX4584);
  nand NAND2_2821(II14934,WX4881,II14933);
  nand NAND2_2822(II14935,WX4584,II14933);
  nand NAND2_2823(II14932,II14934,II14935);
  nand NAND2_2824(II14940,WX4648,II14932);
  nand NAND2_2825(II14941,WX4648,II14940);
  nand NAND2_2826(II14942,II14932,II14940);
  nand NAND2_2827(II14931,II14941,II14942);
  nand NAND2_2828(II14948,WX4712,WX4776);
  nand NAND2_2829(II14949,WX4712,II14948);
  nand NAND2_2830(II14950,WX4776,II14948);
  nand NAND2_2831(II14947,II14949,II14950);
  nand NAND2_2832(II14955,II14931,II14947);
  nand NAND2_2833(II14956,II14931,II14955);
  nand NAND2_2834(II14957,II14947,II14955);
  nand NAND2_2835(WX4809,II14956,II14957);
  nand NAND2_2836(II14964,WX4881,WX4586);
  nand NAND2_2837(II14965,WX4881,II14964);
  nand NAND2_2838(II14966,WX4586,II14964);
  nand NAND2_2839(II14963,II14965,II14966);
  nand NAND2_2840(II14971,WX4650,II14963);
  nand NAND2_2841(II14972,WX4650,II14971);
  nand NAND2_2842(II14973,II14963,II14971);
  nand NAND2_2843(II14962,II14972,II14973);
  nand NAND2_2844(II14979,WX4714,WX4778);
  nand NAND2_2845(II14980,WX4714,II14979);
  nand NAND2_2846(II14981,WX4778,II14979);
  nand NAND2_2847(II14978,II14980,II14981);
  nand NAND2_2848(II14986,II14962,II14978);
  nand NAND2_2849(II14987,II14962,II14986);
  nand NAND2_2850(II14988,II14978,II14986);
  nand NAND2_2851(WX4810,II14987,II14988);
  nand NAND2_2852(II15067,WX4459,WX4364);
  nand NAND2_2853(II15068,WX4459,II15067);
  nand NAND2_2854(II15069,WX4364,II15067);
  nand NAND2_2855(WX4885,II15068,II15069);
  nand NAND2_2856(II15080,WX4460,WX4366);
  nand NAND2_2857(II15081,WX4460,II15080);
  nand NAND2_2858(II15082,WX4366,II15080);
  nand NAND2_2859(WX4892,II15081,II15082);
  nand NAND2_2860(II15093,WX4461,WX4368);
  nand NAND2_2861(II15094,WX4461,II15093);
  nand NAND2_2862(II15095,WX4368,II15093);
  nand NAND2_2863(WX4899,II15094,II15095);
  nand NAND2_2864(II15106,WX4462,WX4370);
  nand NAND2_2865(II15107,WX4462,II15106);
  nand NAND2_2866(II15108,WX4370,II15106);
  nand NAND2_2867(WX4906,II15107,II15108);
  nand NAND2_2868(II15119,WX4463,WX4372);
  nand NAND2_2869(II15120,WX4463,II15119);
  nand NAND2_2870(II15121,WX4372,II15119);
  nand NAND2_2871(WX4913,II15120,II15121);
  nand NAND2_2872(II15132,WX4464,WX4374);
  nand NAND2_2873(II15133,WX4464,II15132);
  nand NAND2_2874(II15134,WX4374,II15132);
  nand NAND2_2875(WX4920,II15133,II15134);
  nand NAND2_2876(II15145,WX4465,WX4376);
  nand NAND2_2877(II15146,WX4465,II15145);
  nand NAND2_2878(II15147,WX4376,II15145);
  nand NAND2_2879(WX4927,II15146,II15147);
  nand NAND2_2880(II15158,WX4466,WX4378);
  nand NAND2_2881(II15159,WX4466,II15158);
  nand NAND2_2882(II15160,WX4378,II15158);
  nand NAND2_2883(WX4934,II15159,II15160);
  nand NAND2_2884(II15171,WX4467,WX4380);
  nand NAND2_2885(II15172,WX4467,II15171);
  nand NAND2_2886(II15173,WX4380,II15171);
  nand NAND2_2887(WX4941,II15172,II15173);
  nand NAND2_2888(II15184,WX4468,WX4382);
  nand NAND2_2889(II15185,WX4468,II15184);
  nand NAND2_2890(II15186,WX4382,II15184);
  nand NAND2_2891(WX4948,II15185,II15186);
  nand NAND2_2892(II15197,WX4469,WX4384);
  nand NAND2_2893(II15198,WX4469,II15197);
  nand NAND2_2894(II15199,WX4384,II15197);
  nand NAND2_2895(WX4955,II15198,II15199);
  nand NAND2_2896(II15210,WX4470,WX4386);
  nand NAND2_2897(II15211,WX4470,II15210);
  nand NAND2_2898(II15212,WX4386,II15210);
  nand NAND2_2899(WX4962,II15211,II15212);
  nand NAND2_2900(II15223,WX4471,WX4388);
  nand NAND2_2901(II15224,WX4471,II15223);
  nand NAND2_2902(II15225,WX4388,II15223);
  nand NAND2_2903(WX4969,II15224,II15225);
  nand NAND2_2904(II15236,WX4472,WX4390);
  nand NAND2_2905(II15237,WX4472,II15236);
  nand NAND2_2906(II15238,WX4390,II15236);
  nand NAND2_2907(WX4976,II15237,II15238);
  nand NAND2_2908(II15249,WX4473,WX4392);
  nand NAND2_2909(II15250,WX4473,II15249);
  nand NAND2_2910(II15251,WX4392,II15249);
  nand NAND2_2911(WX4983,II15250,II15251);
  nand NAND2_2912(II15262,WX4474,WX4394);
  nand NAND2_2913(II15263,WX4474,II15262);
  nand NAND2_2914(II15264,WX4394,II15262);
  nand NAND2_2915(WX4990,II15263,II15264);
  nand NAND2_2916(II15275,WX4475,WX4396);
  nand NAND2_2917(II15276,WX4475,II15275);
  nand NAND2_2918(II15277,WX4396,II15275);
  nand NAND2_2919(WX4997,II15276,II15277);
  nand NAND2_2920(II15288,WX4476,WX4398);
  nand NAND2_2921(II15289,WX4476,II15288);
  nand NAND2_2922(II15290,WX4398,II15288);
  nand NAND2_2923(WX5004,II15289,II15290);
  nand NAND2_2924(II15301,WX4477,WX4400);
  nand NAND2_2925(II15302,WX4477,II15301);
  nand NAND2_2926(II15303,WX4400,II15301);
  nand NAND2_2927(WX5011,II15302,II15303);
  nand NAND2_2928(II15314,WX4478,WX4402);
  nand NAND2_2929(II15315,WX4478,II15314);
  nand NAND2_2930(II15316,WX4402,II15314);
  nand NAND2_2931(WX5018,II15315,II15316);
  nand NAND2_2932(II15327,WX4479,WX4404);
  nand NAND2_2933(II15328,WX4479,II15327);
  nand NAND2_2934(II15329,WX4404,II15327);
  nand NAND2_2935(WX5025,II15328,II15329);
  nand NAND2_2936(II15340,WX4480,WX4406);
  nand NAND2_2937(II15341,WX4480,II15340);
  nand NAND2_2938(II15342,WX4406,II15340);
  nand NAND2_2939(WX5032,II15341,II15342);
  nand NAND2_2940(II15353,WX4481,WX4408);
  nand NAND2_2941(II15354,WX4481,II15353);
  nand NAND2_2942(II15355,WX4408,II15353);
  nand NAND2_2943(WX5039,II15354,II15355);
  nand NAND2_2944(II15366,WX4482,WX4410);
  nand NAND2_2945(II15367,WX4482,II15366);
  nand NAND2_2946(II15368,WX4410,II15366);
  nand NAND2_2947(WX5046,II15367,II15368);
  nand NAND2_2948(II15379,WX4483,WX4412);
  nand NAND2_2949(II15380,WX4483,II15379);
  nand NAND2_2950(II15381,WX4412,II15379);
  nand NAND2_2951(WX5053,II15380,II15381);
  nand NAND2_2952(II15392,WX4484,WX4414);
  nand NAND2_2953(II15393,WX4484,II15392);
  nand NAND2_2954(II15394,WX4414,II15392);
  nand NAND2_2955(WX5060,II15393,II15394);
  nand NAND2_2956(II15405,WX4485,WX4416);
  nand NAND2_2957(II15406,WX4485,II15405);
  nand NAND2_2958(II15407,WX4416,II15405);
  nand NAND2_2959(WX5067,II15406,II15407);
  nand NAND2_2960(II15418,WX4486,WX4418);
  nand NAND2_2961(II15419,WX4486,II15418);
  nand NAND2_2962(II15420,WX4418,II15418);
  nand NAND2_2963(WX5074,II15419,II15420);
  nand NAND2_2964(II15431,WX4487,WX4420);
  nand NAND2_2965(II15432,WX4487,II15431);
  nand NAND2_2966(II15433,WX4420,II15431);
  nand NAND2_2967(WX5081,II15432,II15433);
  nand NAND2_2968(II15444,WX4488,WX4422);
  nand NAND2_2969(II15445,WX4488,II15444);
  nand NAND2_2970(II15446,WX4422,II15444);
  nand NAND2_2971(WX5088,II15445,II15446);
  nand NAND2_2972(II15457,WX4489,WX4424);
  nand NAND2_2973(II15458,WX4489,II15457);
  nand NAND2_2974(II15459,WX4424,II15457);
  nand NAND2_2975(WX5095,II15458,II15459);
  nand NAND2_2976(II15470,WX4490,WX4426);
  nand NAND2_2977(II15471,WX4490,II15470);
  nand NAND2_2978(II15472,WX4426,II15470);
  nand NAND2_2979(WX5102,II15471,II15472);
  nand NAND2_2980(II15485,WX4506,CRC_OUT_6_31);
  nand NAND2_2981(II15486,WX4506,II15485);
  nand NAND2_2982(II15487,CRC_OUT_6_31,II15485);
  nand NAND2_2983(II15484,II15486,II15487);
  nand NAND2_2984(II15492,CRC_OUT_6_15,II15484);
  nand NAND2_2985(II15493,CRC_OUT_6_15,II15492);
  nand NAND2_2986(II15494,II15484,II15492);
  nand NAND2_2987(WX5110,II15493,II15494);
  nand NAND2_2988(II15500,WX4511,CRC_OUT_6_31);
  nand NAND2_2989(II15501,WX4511,II15500);
  nand NAND2_2990(II15502,CRC_OUT_6_31,II15500);
  nand NAND2_2991(II15499,II15501,II15502);
  nand NAND2_2992(II15507,CRC_OUT_6_10,II15499);
  nand NAND2_2993(II15508,CRC_OUT_6_10,II15507);
  nand NAND2_2994(II15509,II15499,II15507);
  nand NAND2_2995(WX5111,II15508,II15509);
  nand NAND2_2996(II15515,WX4518,CRC_OUT_6_31);
  nand NAND2_2997(II15516,WX4518,II15515);
  nand NAND2_2998(II15517,CRC_OUT_6_31,II15515);
  nand NAND2_2999(II15514,II15516,II15517);
  nand NAND2_3000(II15522,CRC_OUT_6_3,II15514);
  nand NAND2_3001(II15523,CRC_OUT_6_3,II15522);
  nand NAND2_3002(II15524,II15514,II15522);
  nand NAND2_3003(WX5112,II15523,II15524);
  nand NAND2_3004(II15529,WX4522,CRC_OUT_6_31);
  nand NAND2_3005(II15530,WX4522,II15529);
  nand NAND2_3006(II15531,CRC_OUT_6_31,II15529);
  nand NAND2_3007(WX5113,II15530,II15531);
  nand NAND2_3008(II15536,WX4491,CRC_OUT_6_30);
  nand NAND2_3009(II15537,WX4491,II15536);
  nand NAND2_3010(II15538,CRC_OUT_6_30,II15536);
  nand NAND2_3011(WX5114,II15537,II15538);
  nand NAND2_3012(II15543,WX4492,CRC_OUT_6_29);
  nand NAND2_3013(II15544,WX4492,II15543);
  nand NAND2_3014(II15545,CRC_OUT_6_29,II15543);
  nand NAND2_3015(WX5115,II15544,II15545);
  nand NAND2_3016(II15550,WX4493,CRC_OUT_6_28);
  nand NAND2_3017(II15551,WX4493,II15550);
  nand NAND2_3018(II15552,CRC_OUT_6_28,II15550);
  nand NAND2_3019(WX5116,II15551,II15552);
  nand NAND2_3020(II15557,WX4494,CRC_OUT_6_27);
  nand NAND2_3021(II15558,WX4494,II15557);
  nand NAND2_3022(II15559,CRC_OUT_6_27,II15557);
  nand NAND2_3023(WX5117,II15558,II15559);
  nand NAND2_3024(II15564,WX4495,CRC_OUT_6_26);
  nand NAND2_3025(II15565,WX4495,II15564);
  nand NAND2_3026(II15566,CRC_OUT_6_26,II15564);
  nand NAND2_3027(WX5118,II15565,II15566);
  nand NAND2_3028(II15571,WX4496,CRC_OUT_6_25);
  nand NAND2_3029(II15572,WX4496,II15571);
  nand NAND2_3030(II15573,CRC_OUT_6_25,II15571);
  nand NAND2_3031(WX5119,II15572,II15573);
  nand NAND2_3032(II15578,WX4497,CRC_OUT_6_24);
  nand NAND2_3033(II15579,WX4497,II15578);
  nand NAND2_3034(II15580,CRC_OUT_6_24,II15578);
  nand NAND2_3035(WX5120,II15579,II15580);
  nand NAND2_3036(II15585,WX4498,CRC_OUT_6_23);
  nand NAND2_3037(II15586,WX4498,II15585);
  nand NAND2_3038(II15587,CRC_OUT_6_23,II15585);
  nand NAND2_3039(WX5121,II15586,II15587);
  nand NAND2_3040(II15592,WX4499,CRC_OUT_6_22);
  nand NAND2_3041(II15593,WX4499,II15592);
  nand NAND2_3042(II15594,CRC_OUT_6_22,II15592);
  nand NAND2_3043(WX5122,II15593,II15594);
  nand NAND2_3044(II15599,WX4500,CRC_OUT_6_21);
  nand NAND2_3045(II15600,WX4500,II15599);
  nand NAND2_3046(II15601,CRC_OUT_6_21,II15599);
  nand NAND2_3047(WX5123,II15600,II15601);
  nand NAND2_3048(II15606,WX4501,CRC_OUT_6_20);
  nand NAND2_3049(II15607,WX4501,II15606);
  nand NAND2_3050(II15608,CRC_OUT_6_20,II15606);
  nand NAND2_3051(WX5124,II15607,II15608);
  nand NAND2_3052(II15613,WX4502,CRC_OUT_6_19);
  nand NAND2_3053(II15614,WX4502,II15613);
  nand NAND2_3054(II15615,CRC_OUT_6_19,II15613);
  nand NAND2_3055(WX5125,II15614,II15615);
  nand NAND2_3056(II15620,WX4503,CRC_OUT_6_18);
  nand NAND2_3057(II15621,WX4503,II15620);
  nand NAND2_3058(II15622,CRC_OUT_6_18,II15620);
  nand NAND2_3059(WX5126,II15621,II15622);
  nand NAND2_3060(II15627,WX4504,CRC_OUT_6_17);
  nand NAND2_3061(II15628,WX4504,II15627);
  nand NAND2_3062(II15629,CRC_OUT_6_17,II15627);
  nand NAND2_3063(WX5127,II15628,II15629);
  nand NAND2_3064(II15634,WX4505,CRC_OUT_6_16);
  nand NAND2_3065(II15635,WX4505,II15634);
  nand NAND2_3066(II15636,CRC_OUT_6_16,II15634);
  nand NAND2_3067(WX5128,II15635,II15636);
  nand NAND2_3068(II15641,WX4507,CRC_OUT_6_14);
  nand NAND2_3069(II15642,WX4507,II15641);
  nand NAND2_3070(II15643,CRC_OUT_6_14,II15641);
  nand NAND2_3071(WX5129,II15642,II15643);
  nand NAND2_3072(II15648,WX4508,CRC_OUT_6_13);
  nand NAND2_3073(II15649,WX4508,II15648);
  nand NAND2_3074(II15650,CRC_OUT_6_13,II15648);
  nand NAND2_3075(WX5130,II15649,II15650);
  nand NAND2_3076(II15655,WX4509,CRC_OUT_6_12);
  nand NAND2_3077(II15656,WX4509,II15655);
  nand NAND2_3078(II15657,CRC_OUT_6_12,II15655);
  nand NAND2_3079(WX5131,II15656,II15657);
  nand NAND2_3080(II15662,WX4510,CRC_OUT_6_11);
  nand NAND2_3081(II15663,WX4510,II15662);
  nand NAND2_3082(II15664,CRC_OUT_6_11,II15662);
  nand NAND2_3083(WX5132,II15663,II15664);
  nand NAND2_3084(II15669,WX4512,CRC_OUT_6_9);
  nand NAND2_3085(II15670,WX4512,II15669);
  nand NAND2_3086(II15671,CRC_OUT_6_9,II15669);
  nand NAND2_3087(WX5133,II15670,II15671);
  nand NAND2_3088(II15676,WX4513,CRC_OUT_6_8);
  nand NAND2_3089(II15677,WX4513,II15676);
  nand NAND2_3090(II15678,CRC_OUT_6_8,II15676);
  nand NAND2_3091(WX5134,II15677,II15678);
  nand NAND2_3092(II15683,WX4514,CRC_OUT_6_7);
  nand NAND2_3093(II15684,WX4514,II15683);
  nand NAND2_3094(II15685,CRC_OUT_6_7,II15683);
  nand NAND2_3095(WX5135,II15684,II15685);
  nand NAND2_3096(II15690,WX4515,CRC_OUT_6_6);
  nand NAND2_3097(II15691,WX4515,II15690);
  nand NAND2_3098(II15692,CRC_OUT_6_6,II15690);
  nand NAND2_3099(WX5136,II15691,II15692);
  nand NAND2_3100(II15697,WX4516,CRC_OUT_6_5);
  nand NAND2_3101(II15698,WX4516,II15697);
  nand NAND2_3102(II15699,CRC_OUT_6_5,II15697);
  nand NAND2_3103(WX5137,II15698,II15699);
  nand NAND2_3104(II15704,WX4517,CRC_OUT_6_4);
  nand NAND2_3105(II15705,WX4517,II15704);
  nand NAND2_3106(II15706,CRC_OUT_6_4,II15704);
  nand NAND2_3107(WX5138,II15705,II15706);
  nand NAND2_3108(II15711,WX4519,CRC_OUT_6_2);
  nand NAND2_3109(II15712,WX4519,II15711);
  nand NAND2_3110(II15713,CRC_OUT_6_2,II15711);
  nand NAND2_3111(WX5139,II15712,II15713);
  nand NAND2_3112(II15718,WX4520,CRC_OUT_6_1);
  nand NAND2_3113(II15719,WX4520,II15718);
  nand NAND2_3114(II15720,CRC_OUT_6_1,II15718);
  nand NAND2_3115(WX5140,II15719,II15720);
  nand NAND2_3116(II15725,WX4521,CRC_OUT_6_0);
  nand NAND2_3117(II15726,WX4521,II15725);
  nand NAND2_3118(II15727,CRC_OUT_6_0,II15725);
  nand NAND2_3119(WX5141,II15726,II15727);
  nand NAND2_3120(II18008,WX6173,WX5817);
  nand NAND2_3121(II18009,WX6173,II18008);
  nand NAND2_3122(II18010,WX5817,II18008);
  nand NAND2_3123(II18007,II18009,II18010);
  nand NAND2_3124(II18015,WX5881,II18007);
  nand NAND2_3125(II18016,WX5881,II18015);
  nand NAND2_3126(II18017,II18007,II18015);
  nand NAND2_3127(II18006,II18016,II18017);
  nand NAND2_3128(II18023,WX5945,WX6009);
  nand NAND2_3129(II18024,WX5945,II18023);
  nand NAND2_3130(II18025,WX6009,II18023);
  nand NAND2_3131(II18022,II18024,II18025);
  nand NAND2_3132(II18030,II18006,II18022);
  nand NAND2_3133(II18031,II18006,II18030);
  nand NAND2_3134(II18032,II18022,II18030);
  nand NAND2_3135(WX6072,II18031,II18032);
  nand NAND2_3136(II18039,WX6173,WX5819);
  nand NAND2_3137(II18040,WX6173,II18039);
  nand NAND2_3138(II18041,WX5819,II18039);
  nand NAND2_3139(II18038,II18040,II18041);
  nand NAND2_3140(II18046,WX5883,II18038);
  nand NAND2_3141(II18047,WX5883,II18046);
  nand NAND2_3142(II18048,II18038,II18046);
  nand NAND2_3143(II18037,II18047,II18048);
  nand NAND2_3144(II18054,WX5947,WX6011);
  nand NAND2_3145(II18055,WX5947,II18054);
  nand NAND2_3146(II18056,WX6011,II18054);
  nand NAND2_3147(II18053,II18055,II18056);
  nand NAND2_3148(II18061,II18037,II18053);
  nand NAND2_3149(II18062,II18037,II18061);
  nand NAND2_3150(II18063,II18053,II18061);
  nand NAND2_3151(WX6073,II18062,II18063);
  nand NAND2_3152(II18070,WX6173,WX5821);
  nand NAND2_3153(II18071,WX6173,II18070);
  nand NAND2_3154(II18072,WX5821,II18070);
  nand NAND2_3155(II18069,II18071,II18072);
  nand NAND2_3156(II18077,WX5885,II18069);
  nand NAND2_3157(II18078,WX5885,II18077);
  nand NAND2_3158(II18079,II18069,II18077);
  nand NAND2_3159(II18068,II18078,II18079);
  nand NAND2_3160(II18085,WX5949,WX6013);
  nand NAND2_3161(II18086,WX5949,II18085);
  nand NAND2_3162(II18087,WX6013,II18085);
  nand NAND2_3163(II18084,II18086,II18087);
  nand NAND2_3164(II18092,II18068,II18084);
  nand NAND2_3165(II18093,II18068,II18092);
  nand NAND2_3166(II18094,II18084,II18092);
  nand NAND2_3167(WX6074,II18093,II18094);
  nand NAND2_3168(II18101,WX6173,WX5823);
  nand NAND2_3169(II18102,WX6173,II18101);
  nand NAND2_3170(II18103,WX5823,II18101);
  nand NAND2_3171(II18100,II18102,II18103);
  nand NAND2_3172(II18108,WX5887,II18100);
  nand NAND2_3173(II18109,WX5887,II18108);
  nand NAND2_3174(II18110,II18100,II18108);
  nand NAND2_3175(II18099,II18109,II18110);
  nand NAND2_3176(II18116,WX5951,WX6015);
  nand NAND2_3177(II18117,WX5951,II18116);
  nand NAND2_3178(II18118,WX6015,II18116);
  nand NAND2_3179(II18115,II18117,II18118);
  nand NAND2_3180(II18123,II18099,II18115);
  nand NAND2_3181(II18124,II18099,II18123);
  nand NAND2_3182(II18125,II18115,II18123);
  nand NAND2_3183(WX6075,II18124,II18125);
  nand NAND2_3184(II18132,WX6173,WX5825);
  nand NAND2_3185(II18133,WX6173,II18132);
  nand NAND2_3186(II18134,WX5825,II18132);
  nand NAND2_3187(II18131,II18133,II18134);
  nand NAND2_3188(II18139,WX5889,II18131);
  nand NAND2_3189(II18140,WX5889,II18139);
  nand NAND2_3190(II18141,II18131,II18139);
  nand NAND2_3191(II18130,II18140,II18141);
  nand NAND2_3192(II18147,WX5953,WX6017);
  nand NAND2_3193(II18148,WX5953,II18147);
  nand NAND2_3194(II18149,WX6017,II18147);
  nand NAND2_3195(II18146,II18148,II18149);
  nand NAND2_3196(II18154,II18130,II18146);
  nand NAND2_3197(II18155,II18130,II18154);
  nand NAND2_3198(II18156,II18146,II18154);
  nand NAND2_3199(WX6076,II18155,II18156);
  nand NAND2_3200(II18163,WX6173,WX5827);
  nand NAND2_3201(II18164,WX6173,II18163);
  nand NAND2_3202(II18165,WX5827,II18163);
  nand NAND2_3203(II18162,II18164,II18165);
  nand NAND2_3204(II18170,WX5891,II18162);
  nand NAND2_3205(II18171,WX5891,II18170);
  nand NAND2_3206(II18172,II18162,II18170);
  nand NAND2_3207(II18161,II18171,II18172);
  nand NAND2_3208(II18178,WX5955,WX6019);
  nand NAND2_3209(II18179,WX5955,II18178);
  nand NAND2_3210(II18180,WX6019,II18178);
  nand NAND2_3211(II18177,II18179,II18180);
  nand NAND2_3212(II18185,II18161,II18177);
  nand NAND2_3213(II18186,II18161,II18185);
  nand NAND2_3214(II18187,II18177,II18185);
  nand NAND2_3215(WX6077,II18186,II18187);
  nand NAND2_3216(II18194,WX6173,WX5829);
  nand NAND2_3217(II18195,WX6173,II18194);
  nand NAND2_3218(II18196,WX5829,II18194);
  nand NAND2_3219(II18193,II18195,II18196);
  nand NAND2_3220(II18201,WX5893,II18193);
  nand NAND2_3221(II18202,WX5893,II18201);
  nand NAND2_3222(II18203,II18193,II18201);
  nand NAND2_3223(II18192,II18202,II18203);
  nand NAND2_3224(II18209,WX5957,WX6021);
  nand NAND2_3225(II18210,WX5957,II18209);
  nand NAND2_3226(II18211,WX6021,II18209);
  nand NAND2_3227(II18208,II18210,II18211);
  nand NAND2_3228(II18216,II18192,II18208);
  nand NAND2_3229(II18217,II18192,II18216);
  nand NAND2_3230(II18218,II18208,II18216);
  nand NAND2_3231(WX6078,II18217,II18218);
  nand NAND2_3232(II18225,WX6173,WX5831);
  nand NAND2_3233(II18226,WX6173,II18225);
  nand NAND2_3234(II18227,WX5831,II18225);
  nand NAND2_3235(II18224,II18226,II18227);
  nand NAND2_3236(II18232,WX5895,II18224);
  nand NAND2_3237(II18233,WX5895,II18232);
  nand NAND2_3238(II18234,II18224,II18232);
  nand NAND2_3239(II18223,II18233,II18234);
  nand NAND2_3240(II18240,WX5959,WX6023);
  nand NAND2_3241(II18241,WX5959,II18240);
  nand NAND2_3242(II18242,WX6023,II18240);
  nand NAND2_3243(II18239,II18241,II18242);
  nand NAND2_3244(II18247,II18223,II18239);
  nand NAND2_3245(II18248,II18223,II18247);
  nand NAND2_3246(II18249,II18239,II18247);
  nand NAND2_3247(WX6079,II18248,II18249);
  nand NAND2_3248(II18256,WX6173,WX5833);
  nand NAND2_3249(II18257,WX6173,II18256);
  nand NAND2_3250(II18258,WX5833,II18256);
  nand NAND2_3251(II18255,II18257,II18258);
  nand NAND2_3252(II18263,WX5897,II18255);
  nand NAND2_3253(II18264,WX5897,II18263);
  nand NAND2_3254(II18265,II18255,II18263);
  nand NAND2_3255(II18254,II18264,II18265);
  nand NAND2_3256(II18271,WX5961,WX6025);
  nand NAND2_3257(II18272,WX5961,II18271);
  nand NAND2_3258(II18273,WX6025,II18271);
  nand NAND2_3259(II18270,II18272,II18273);
  nand NAND2_3260(II18278,II18254,II18270);
  nand NAND2_3261(II18279,II18254,II18278);
  nand NAND2_3262(II18280,II18270,II18278);
  nand NAND2_3263(WX6080,II18279,II18280);
  nand NAND2_3264(II18287,WX6173,WX5835);
  nand NAND2_3265(II18288,WX6173,II18287);
  nand NAND2_3266(II18289,WX5835,II18287);
  nand NAND2_3267(II18286,II18288,II18289);
  nand NAND2_3268(II18294,WX5899,II18286);
  nand NAND2_3269(II18295,WX5899,II18294);
  nand NAND2_3270(II18296,II18286,II18294);
  nand NAND2_3271(II18285,II18295,II18296);
  nand NAND2_3272(II18302,WX5963,WX6027);
  nand NAND2_3273(II18303,WX5963,II18302);
  nand NAND2_3274(II18304,WX6027,II18302);
  nand NAND2_3275(II18301,II18303,II18304);
  nand NAND2_3276(II18309,II18285,II18301);
  nand NAND2_3277(II18310,II18285,II18309);
  nand NAND2_3278(II18311,II18301,II18309);
  nand NAND2_3279(WX6081,II18310,II18311);
  nand NAND2_3280(II18318,WX6173,WX5837);
  nand NAND2_3281(II18319,WX6173,II18318);
  nand NAND2_3282(II18320,WX5837,II18318);
  nand NAND2_3283(II18317,II18319,II18320);
  nand NAND2_3284(II18325,WX5901,II18317);
  nand NAND2_3285(II18326,WX5901,II18325);
  nand NAND2_3286(II18327,II18317,II18325);
  nand NAND2_3287(II18316,II18326,II18327);
  nand NAND2_3288(II18333,WX5965,WX6029);
  nand NAND2_3289(II18334,WX5965,II18333);
  nand NAND2_3290(II18335,WX6029,II18333);
  nand NAND2_3291(II18332,II18334,II18335);
  nand NAND2_3292(II18340,II18316,II18332);
  nand NAND2_3293(II18341,II18316,II18340);
  nand NAND2_3294(II18342,II18332,II18340);
  nand NAND2_3295(WX6082,II18341,II18342);
  nand NAND2_3296(II18349,WX6173,WX5839);
  nand NAND2_3297(II18350,WX6173,II18349);
  nand NAND2_3298(II18351,WX5839,II18349);
  nand NAND2_3299(II18348,II18350,II18351);
  nand NAND2_3300(II18356,WX5903,II18348);
  nand NAND2_3301(II18357,WX5903,II18356);
  nand NAND2_3302(II18358,II18348,II18356);
  nand NAND2_3303(II18347,II18357,II18358);
  nand NAND2_3304(II18364,WX5967,WX6031);
  nand NAND2_3305(II18365,WX5967,II18364);
  nand NAND2_3306(II18366,WX6031,II18364);
  nand NAND2_3307(II18363,II18365,II18366);
  nand NAND2_3308(II18371,II18347,II18363);
  nand NAND2_3309(II18372,II18347,II18371);
  nand NAND2_3310(II18373,II18363,II18371);
  nand NAND2_3311(WX6083,II18372,II18373);
  nand NAND2_3312(II18380,WX6173,WX5841);
  nand NAND2_3313(II18381,WX6173,II18380);
  nand NAND2_3314(II18382,WX5841,II18380);
  nand NAND2_3315(II18379,II18381,II18382);
  nand NAND2_3316(II18387,WX5905,II18379);
  nand NAND2_3317(II18388,WX5905,II18387);
  nand NAND2_3318(II18389,II18379,II18387);
  nand NAND2_3319(II18378,II18388,II18389);
  nand NAND2_3320(II18395,WX5969,WX6033);
  nand NAND2_3321(II18396,WX5969,II18395);
  nand NAND2_3322(II18397,WX6033,II18395);
  nand NAND2_3323(II18394,II18396,II18397);
  nand NAND2_3324(II18402,II18378,II18394);
  nand NAND2_3325(II18403,II18378,II18402);
  nand NAND2_3326(II18404,II18394,II18402);
  nand NAND2_3327(WX6084,II18403,II18404);
  nand NAND2_3328(II18411,WX6173,WX5843);
  nand NAND2_3329(II18412,WX6173,II18411);
  nand NAND2_3330(II18413,WX5843,II18411);
  nand NAND2_3331(II18410,II18412,II18413);
  nand NAND2_3332(II18418,WX5907,II18410);
  nand NAND2_3333(II18419,WX5907,II18418);
  nand NAND2_3334(II18420,II18410,II18418);
  nand NAND2_3335(II18409,II18419,II18420);
  nand NAND2_3336(II18426,WX5971,WX6035);
  nand NAND2_3337(II18427,WX5971,II18426);
  nand NAND2_3338(II18428,WX6035,II18426);
  nand NAND2_3339(II18425,II18427,II18428);
  nand NAND2_3340(II18433,II18409,II18425);
  nand NAND2_3341(II18434,II18409,II18433);
  nand NAND2_3342(II18435,II18425,II18433);
  nand NAND2_3343(WX6085,II18434,II18435);
  nand NAND2_3344(II18442,WX6173,WX5845);
  nand NAND2_3345(II18443,WX6173,II18442);
  nand NAND2_3346(II18444,WX5845,II18442);
  nand NAND2_3347(II18441,II18443,II18444);
  nand NAND2_3348(II18449,WX5909,II18441);
  nand NAND2_3349(II18450,WX5909,II18449);
  nand NAND2_3350(II18451,II18441,II18449);
  nand NAND2_3351(II18440,II18450,II18451);
  nand NAND2_3352(II18457,WX5973,WX6037);
  nand NAND2_3353(II18458,WX5973,II18457);
  nand NAND2_3354(II18459,WX6037,II18457);
  nand NAND2_3355(II18456,II18458,II18459);
  nand NAND2_3356(II18464,II18440,II18456);
  nand NAND2_3357(II18465,II18440,II18464);
  nand NAND2_3358(II18466,II18456,II18464);
  nand NAND2_3359(WX6086,II18465,II18466);
  nand NAND2_3360(II18473,WX6173,WX5847);
  nand NAND2_3361(II18474,WX6173,II18473);
  nand NAND2_3362(II18475,WX5847,II18473);
  nand NAND2_3363(II18472,II18474,II18475);
  nand NAND2_3364(II18480,WX5911,II18472);
  nand NAND2_3365(II18481,WX5911,II18480);
  nand NAND2_3366(II18482,II18472,II18480);
  nand NAND2_3367(II18471,II18481,II18482);
  nand NAND2_3368(II18488,WX5975,WX6039);
  nand NAND2_3369(II18489,WX5975,II18488);
  nand NAND2_3370(II18490,WX6039,II18488);
  nand NAND2_3371(II18487,II18489,II18490);
  nand NAND2_3372(II18495,II18471,II18487);
  nand NAND2_3373(II18496,II18471,II18495);
  nand NAND2_3374(II18497,II18487,II18495);
  nand NAND2_3375(WX6087,II18496,II18497);
  nand NAND2_3376(II18504,WX6174,WX5849);
  nand NAND2_3377(II18505,WX6174,II18504);
  nand NAND2_3378(II18506,WX5849,II18504);
  nand NAND2_3379(II18503,II18505,II18506);
  nand NAND2_3380(II18511,WX5913,II18503);
  nand NAND2_3381(II18512,WX5913,II18511);
  nand NAND2_3382(II18513,II18503,II18511);
  nand NAND2_3383(II18502,II18512,II18513);
  nand NAND2_3384(II18519,WX5977,WX6041);
  nand NAND2_3385(II18520,WX5977,II18519);
  nand NAND2_3386(II18521,WX6041,II18519);
  nand NAND2_3387(II18518,II18520,II18521);
  nand NAND2_3388(II18526,II18502,II18518);
  nand NAND2_3389(II18527,II18502,II18526);
  nand NAND2_3390(II18528,II18518,II18526);
  nand NAND2_3391(WX6088,II18527,II18528);
  nand NAND2_3392(II18535,WX6174,WX5851);
  nand NAND2_3393(II18536,WX6174,II18535);
  nand NAND2_3394(II18537,WX5851,II18535);
  nand NAND2_3395(II18534,II18536,II18537);
  nand NAND2_3396(II18542,WX5915,II18534);
  nand NAND2_3397(II18543,WX5915,II18542);
  nand NAND2_3398(II18544,II18534,II18542);
  nand NAND2_3399(II18533,II18543,II18544);
  nand NAND2_3400(II18550,WX5979,WX6043);
  nand NAND2_3401(II18551,WX5979,II18550);
  nand NAND2_3402(II18552,WX6043,II18550);
  nand NAND2_3403(II18549,II18551,II18552);
  nand NAND2_3404(II18557,II18533,II18549);
  nand NAND2_3405(II18558,II18533,II18557);
  nand NAND2_3406(II18559,II18549,II18557);
  nand NAND2_3407(WX6089,II18558,II18559);
  nand NAND2_3408(II18566,WX6174,WX5853);
  nand NAND2_3409(II18567,WX6174,II18566);
  nand NAND2_3410(II18568,WX5853,II18566);
  nand NAND2_3411(II18565,II18567,II18568);
  nand NAND2_3412(II18573,WX5917,II18565);
  nand NAND2_3413(II18574,WX5917,II18573);
  nand NAND2_3414(II18575,II18565,II18573);
  nand NAND2_3415(II18564,II18574,II18575);
  nand NAND2_3416(II18581,WX5981,WX6045);
  nand NAND2_3417(II18582,WX5981,II18581);
  nand NAND2_3418(II18583,WX6045,II18581);
  nand NAND2_3419(II18580,II18582,II18583);
  nand NAND2_3420(II18588,II18564,II18580);
  nand NAND2_3421(II18589,II18564,II18588);
  nand NAND2_3422(II18590,II18580,II18588);
  nand NAND2_3423(WX6090,II18589,II18590);
  nand NAND2_3424(II18597,WX6174,WX5855);
  nand NAND2_3425(II18598,WX6174,II18597);
  nand NAND2_3426(II18599,WX5855,II18597);
  nand NAND2_3427(II18596,II18598,II18599);
  nand NAND2_3428(II18604,WX5919,II18596);
  nand NAND2_3429(II18605,WX5919,II18604);
  nand NAND2_3430(II18606,II18596,II18604);
  nand NAND2_3431(II18595,II18605,II18606);
  nand NAND2_3432(II18612,WX5983,WX6047);
  nand NAND2_3433(II18613,WX5983,II18612);
  nand NAND2_3434(II18614,WX6047,II18612);
  nand NAND2_3435(II18611,II18613,II18614);
  nand NAND2_3436(II18619,II18595,II18611);
  nand NAND2_3437(II18620,II18595,II18619);
  nand NAND2_3438(II18621,II18611,II18619);
  nand NAND2_3439(WX6091,II18620,II18621);
  nand NAND2_3440(II18628,WX6174,WX5857);
  nand NAND2_3441(II18629,WX6174,II18628);
  nand NAND2_3442(II18630,WX5857,II18628);
  nand NAND2_3443(II18627,II18629,II18630);
  nand NAND2_3444(II18635,WX5921,II18627);
  nand NAND2_3445(II18636,WX5921,II18635);
  nand NAND2_3446(II18637,II18627,II18635);
  nand NAND2_3447(II18626,II18636,II18637);
  nand NAND2_3448(II18643,WX5985,WX6049);
  nand NAND2_3449(II18644,WX5985,II18643);
  nand NAND2_3450(II18645,WX6049,II18643);
  nand NAND2_3451(II18642,II18644,II18645);
  nand NAND2_3452(II18650,II18626,II18642);
  nand NAND2_3453(II18651,II18626,II18650);
  nand NAND2_3454(II18652,II18642,II18650);
  nand NAND2_3455(WX6092,II18651,II18652);
  nand NAND2_3456(II18659,WX6174,WX5859);
  nand NAND2_3457(II18660,WX6174,II18659);
  nand NAND2_3458(II18661,WX5859,II18659);
  nand NAND2_3459(II18658,II18660,II18661);
  nand NAND2_3460(II18666,WX5923,II18658);
  nand NAND2_3461(II18667,WX5923,II18666);
  nand NAND2_3462(II18668,II18658,II18666);
  nand NAND2_3463(II18657,II18667,II18668);
  nand NAND2_3464(II18674,WX5987,WX6051);
  nand NAND2_3465(II18675,WX5987,II18674);
  nand NAND2_3466(II18676,WX6051,II18674);
  nand NAND2_3467(II18673,II18675,II18676);
  nand NAND2_3468(II18681,II18657,II18673);
  nand NAND2_3469(II18682,II18657,II18681);
  nand NAND2_3470(II18683,II18673,II18681);
  nand NAND2_3471(WX6093,II18682,II18683);
  nand NAND2_3472(II18690,WX6174,WX5861);
  nand NAND2_3473(II18691,WX6174,II18690);
  nand NAND2_3474(II18692,WX5861,II18690);
  nand NAND2_3475(II18689,II18691,II18692);
  nand NAND2_3476(II18697,WX5925,II18689);
  nand NAND2_3477(II18698,WX5925,II18697);
  nand NAND2_3478(II18699,II18689,II18697);
  nand NAND2_3479(II18688,II18698,II18699);
  nand NAND2_3480(II18705,WX5989,WX6053);
  nand NAND2_3481(II18706,WX5989,II18705);
  nand NAND2_3482(II18707,WX6053,II18705);
  nand NAND2_3483(II18704,II18706,II18707);
  nand NAND2_3484(II18712,II18688,II18704);
  nand NAND2_3485(II18713,II18688,II18712);
  nand NAND2_3486(II18714,II18704,II18712);
  nand NAND2_3487(WX6094,II18713,II18714);
  nand NAND2_3488(II18721,WX6174,WX5863);
  nand NAND2_3489(II18722,WX6174,II18721);
  nand NAND2_3490(II18723,WX5863,II18721);
  nand NAND2_3491(II18720,II18722,II18723);
  nand NAND2_3492(II18728,WX5927,II18720);
  nand NAND2_3493(II18729,WX5927,II18728);
  nand NAND2_3494(II18730,II18720,II18728);
  nand NAND2_3495(II18719,II18729,II18730);
  nand NAND2_3496(II18736,WX5991,WX6055);
  nand NAND2_3497(II18737,WX5991,II18736);
  nand NAND2_3498(II18738,WX6055,II18736);
  nand NAND2_3499(II18735,II18737,II18738);
  nand NAND2_3500(II18743,II18719,II18735);
  nand NAND2_3501(II18744,II18719,II18743);
  nand NAND2_3502(II18745,II18735,II18743);
  nand NAND2_3503(WX6095,II18744,II18745);
  nand NAND2_3504(II18752,WX6174,WX5865);
  nand NAND2_3505(II18753,WX6174,II18752);
  nand NAND2_3506(II18754,WX5865,II18752);
  nand NAND2_3507(II18751,II18753,II18754);
  nand NAND2_3508(II18759,WX5929,II18751);
  nand NAND2_3509(II18760,WX5929,II18759);
  nand NAND2_3510(II18761,II18751,II18759);
  nand NAND2_3511(II18750,II18760,II18761);
  nand NAND2_3512(II18767,WX5993,WX6057);
  nand NAND2_3513(II18768,WX5993,II18767);
  nand NAND2_3514(II18769,WX6057,II18767);
  nand NAND2_3515(II18766,II18768,II18769);
  nand NAND2_3516(II18774,II18750,II18766);
  nand NAND2_3517(II18775,II18750,II18774);
  nand NAND2_3518(II18776,II18766,II18774);
  nand NAND2_3519(WX6096,II18775,II18776);
  nand NAND2_3520(II18783,WX6174,WX5867);
  nand NAND2_3521(II18784,WX6174,II18783);
  nand NAND2_3522(II18785,WX5867,II18783);
  nand NAND2_3523(II18782,II18784,II18785);
  nand NAND2_3524(II18790,WX5931,II18782);
  nand NAND2_3525(II18791,WX5931,II18790);
  nand NAND2_3526(II18792,II18782,II18790);
  nand NAND2_3527(II18781,II18791,II18792);
  nand NAND2_3528(II18798,WX5995,WX6059);
  nand NAND2_3529(II18799,WX5995,II18798);
  nand NAND2_3530(II18800,WX6059,II18798);
  nand NAND2_3531(II18797,II18799,II18800);
  nand NAND2_3532(II18805,II18781,II18797);
  nand NAND2_3533(II18806,II18781,II18805);
  nand NAND2_3534(II18807,II18797,II18805);
  nand NAND2_3535(WX6097,II18806,II18807);
  nand NAND2_3536(II18814,WX6174,WX5869);
  nand NAND2_3537(II18815,WX6174,II18814);
  nand NAND2_3538(II18816,WX5869,II18814);
  nand NAND2_3539(II18813,II18815,II18816);
  nand NAND2_3540(II18821,WX5933,II18813);
  nand NAND2_3541(II18822,WX5933,II18821);
  nand NAND2_3542(II18823,II18813,II18821);
  nand NAND2_3543(II18812,II18822,II18823);
  nand NAND2_3544(II18829,WX5997,WX6061);
  nand NAND2_3545(II18830,WX5997,II18829);
  nand NAND2_3546(II18831,WX6061,II18829);
  nand NAND2_3547(II18828,II18830,II18831);
  nand NAND2_3548(II18836,II18812,II18828);
  nand NAND2_3549(II18837,II18812,II18836);
  nand NAND2_3550(II18838,II18828,II18836);
  nand NAND2_3551(WX6098,II18837,II18838);
  nand NAND2_3552(II18845,WX6174,WX5871);
  nand NAND2_3553(II18846,WX6174,II18845);
  nand NAND2_3554(II18847,WX5871,II18845);
  nand NAND2_3555(II18844,II18846,II18847);
  nand NAND2_3556(II18852,WX5935,II18844);
  nand NAND2_3557(II18853,WX5935,II18852);
  nand NAND2_3558(II18854,II18844,II18852);
  nand NAND2_3559(II18843,II18853,II18854);
  nand NAND2_3560(II18860,WX5999,WX6063);
  nand NAND2_3561(II18861,WX5999,II18860);
  nand NAND2_3562(II18862,WX6063,II18860);
  nand NAND2_3563(II18859,II18861,II18862);
  nand NAND2_3564(II18867,II18843,II18859);
  nand NAND2_3565(II18868,II18843,II18867);
  nand NAND2_3566(II18869,II18859,II18867);
  nand NAND2_3567(WX6099,II18868,II18869);
  nand NAND2_3568(II18876,WX6174,WX5873);
  nand NAND2_3569(II18877,WX6174,II18876);
  nand NAND2_3570(II18878,WX5873,II18876);
  nand NAND2_3571(II18875,II18877,II18878);
  nand NAND2_3572(II18883,WX5937,II18875);
  nand NAND2_3573(II18884,WX5937,II18883);
  nand NAND2_3574(II18885,II18875,II18883);
  nand NAND2_3575(II18874,II18884,II18885);
  nand NAND2_3576(II18891,WX6001,WX6065);
  nand NAND2_3577(II18892,WX6001,II18891);
  nand NAND2_3578(II18893,WX6065,II18891);
  nand NAND2_3579(II18890,II18892,II18893);
  nand NAND2_3580(II18898,II18874,II18890);
  nand NAND2_3581(II18899,II18874,II18898);
  nand NAND2_3582(II18900,II18890,II18898);
  nand NAND2_3583(WX6100,II18899,II18900);
  nand NAND2_3584(II18907,WX6174,WX5875);
  nand NAND2_3585(II18908,WX6174,II18907);
  nand NAND2_3586(II18909,WX5875,II18907);
  nand NAND2_3587(II18906,II18908,II18909);
  nand NAND2_3588(II18914,WX5939,II18906);
  nand NAND2_3589(II18915,WX5939,II18914);
  nand NAND2_3590(II18916,II18906,II18914);
  nand NAND2_3591(II18905,II18915,II18916);
  nand NAND2_3592(II18922,WX6003,WX6067);
  nand NAND2_3593(II18923,WX6003,II18922);
  nand NAND2_3594(II18924,WX6067,II18922);
  nand NAND2_3595(II18921,II18923,II18924);
  nand NAND2_3596(II18929,II18905,II18921);
  nand NAND2_3597(II18930,II18905,II18929);
  nand NAND2_3598(II18931,II18921,II18929);
  nand NAND2_3599(WX6101,II18930,II18931);
  nand NAND2_3600(II18938,WX6174,WX5877);
  nand NAND2_3601(II18939,WX6174,II18938);
  nand NAND2_3602(II18940,WX5877,II18938);
  nand NAND2_3603(II18937,II18939,II18940);
  nand NAND2_3604(II18945,WX5941,II18937);
  nand NAND2_3605(II18946,WX5941,II18945);
  nand NAND2_3606(II18947,II18937,II18945);
  nand NAND2_3607(II18936,II18946,II18947);
  nand NAND2_3608(II18953,WX6005,WX6069);
  nand NAND2_3609(II18954,WX6005,II18953);
  nand NAND2_3610(II18955,WX6069,II18953);
  nand NAND2_3611(II18952,II18954,II18955);
  nand NAND2_3612(II18960,II18936,II18952);
  nand NAND2_3613(II18961,II18936,II18960);
  nand NAND2_3614(II18962,II18952,II18960);
  nand NAND2_3615(WX6102,II18961,II18962);
  nand NAND2_3616(II18969,WX6174,WX5879);
  nand NAND2_3617(II18970,WX6174,II18969);
  nand NAND2_3618(II18971,WX5879,II18969);
  nand NAND2_3619(II18968,II18970,II18971);
  nand NAND2_3620(II18976,WX5943,II18968);
  nand NAND2_3621(II18977,WX5943,II18976);
  nand NAND2_3622(II18978,II18968,II18976);
  nand NAND2_3623(II18967,II18977,II18978);
  nand NAND2_3624(II18984,WX6007,WX6071);
  nand NAND2_3625(II18985,WX6007,II18984);
  nand NAND2_3626(II18986,WX6071,II18984);
  nand NAND2_3627(II18983,II18985,II18986);
  nand NAND2_3628(II18991,II18967,II18983);
  nand NAND2_3629(II18992,II18967,II18991);
  nand NAND2_3630(II18993,II18983,II18991);
  nand NAND2_3631(WX6103,II18992,II18993);
  nand NAND2_3632(II19072,WX5752,WX5657);
  nand NAND2_3633(II19073,WX5752,II19072);
  nand NAND2_3634(II19074,WX5657,II19072);
  nand NAND2_3635(WX6178,II19073,II19074);
  nand NAND2_3636(II19085,WX5753,WX5659);
  nand NAND2_3637(II19086,WX5753,II19085);
  nand NAND2_3638(II19087,WX5659,II19085);
  nand NAND2_3639(WX6185,II19086,II19087);
  nand NAND2_3640(II19098,WX5754,WX5661);
  nand NAND2_3641(II19099,WX5754,II19098);
  nand NAND2_3642(II19100,WX5661,II19098);
  nand NAND2_3643(WX6192,II19099,II19100);
  nand NAND2_3644(II19111,WX5755,WX5663);
  nand NAND2_3645(II19112,WX5755,II19111);
  nand NAND2_3646(II19113,WX5663,II19111);
  nand NAND2_3647(WX6199,II19112,II19113);
  nand NAND2_3648(II19124,WX5756,WX5665);
  nand NAND2_3649(II19125,WX5756,II19124);
  nand NAND2_3650(II19126,WX5665,II19124);
  nand NAND2_3651(WX6206,II19125,II19126);
  nand NAND2_3652(II19137,WX5757,WX5667);
  nand NAND2_3653(II19138,WX5757,II19137);
  nand NAND2_3654(II19139,WX5667,II19137);
  nand NAND2_3655(WX6213,II19138,II19139);
  nand NAND2_3656(II19150,WX5758,WX5669);
  nand NAND2_3657(II19151,WX5758,II19150);
  nand NAND2_3658(II19152,WX5669,II19150);
  nand NAND2_3659(WX6220,II19151,II19152);
  nand NAND2_3660(II19163,WX5759,WX5671);
  nand NAND2_3661(II19164,WX5759,II19163);
  nand NAND2_3662(II19165,WX5671,II19163);
  nand NAND2_3663(WX6227,II19164,II19165);
  nand NAND2_3664(II19176,WX5760,WX5673);
  nand NAND2_3665(II19177,WX5760,II19176);
  nand NAND2_3666(II19178,WX5673,II19176);
  nand NAND2_3667(WX6234,II19177,II19178);
  nand NAND2_3668(II19189,WX5761,WX5675);
  nand NAND2_3669(II19190,WX5761,II19189);
  nand NAND2_3670(II19191,WX5675,II19189);
  nand NAND2_3671(WX6241,II19190,II19191);
  nand NAND2_3672(II19202,WX5762,WX5677);
  nand NAND2_3673(II19203,WX5762,II19202);
  nand NAND2_3674(II19204,WX5677,II19202);
  nand NAND2_3675(WX6248,II19203,II19204);
  nand NAND2_3676(II19215,WX5763,WX5679);
  nand NAND2_3677(II19216,WX5763,II19215);
  nand NAND2_3678(II19217,WX5679,II19215);
  nand NAND2_3679(WX6255,II19216,II19217);
  nand NAND2_3680(II19228,WX5764,WX5681);
  nand NAND2_3681(II19229,WX5764,II19228);
  nand NAND2_3682(II19230,WX5681,II19228);
  nand NAND2_3683(WX6262,II19229,II19230);
  nand NAND2_3684(II19241,WX5765,WX5683);
  nand NAND2_3685(II19242,WX5765,II19241);
  nand NAND2_3686(II19243,WX5683,II19241);
  nand NAND2_3687(WX6269,II19242,II19243);
  nand NAND2_3688(II19254,WX5766,WX5685);
  nand NAND2_3689(II19255,WX5766,II19254);
  nand NAND2_3690(II19256,WX5685,II19254);
  nand NAND2_3691(WX6276,II19255,II19256);
  nand NAND2_3692(II19267,WX5767,WX5687);
  nand NAND2_3693(II19268,WX5767,II19267);
  nand NAND2_3694(II19269,WX5687,II19267);
  nand NAND2_3695(WX6283,II19268,II19269);
  nand NAND2_3696(II19280,WX5768,WX5689);
  nand NAND2_3697(II19281,WX5768,II19280);
  nand NAND2_3698(II19282,WX5689,II19280);
  nand NAND2_3699(WX6290,II19281,II19282);
  nand NAND2_3700(II19293,WX5769,WX5691);
  nand NAND2_3701(II19294,WX5769,II19293);
  nand NAND2_3702(II19295,WX5691,II19293);
  nand NAND2_3703(WX6297,II19294,II19295);
  nand NAND2_3704(II19306,WX5770,WX5693);
  nand NAND2_3705(II19307,WX5770,II19306);
  nand NAND2_3706(II19308,WX5693,II19306);
  nand NAND2_3707(WX6304,II19307,II19308);
  nand NAND2_3708(II19319,WX5771,WX5695);
  nand NAND2_3709(II19320,WX5771,II19319);
  nand NAND2_3710(II19321,WX5695,II19319);
  nand NAND2_3711(WX6311,II19320,II19321);
  nand NAND2_3712(II19332,WX5772,WX5697);
  nand NAND2_3713(II19333,WX5772,II19332);
  nand NAND2_3714(II19334,WX5697,II19332);
  nand NAND2_3715(WX6318,II19333,II19334);
  nand NAND2_3716(II19345,WX5773,WX5699);
  nand NAND2_3717(II19346,WX5773,II19345);
  nand NAND2_3718(II19347,WX5699,II19345);
  nand NAND2_3719(WX6325,II19346,II19347);
  nand NAND2_3720(II19358,WX5774,WX5701);
  nand NAND2_3721(II19359,WX5774,II19358);
  nand NAND2_3722(II19360,WX5701,II19358);
  nand NAND2_3723(WX6332,II19359,II19360);
  nand NAND2_3724(II19371,WX5775,WX5703);
  nand NAND2_3725(II19372,WX5775,II19371);
  nand NAND2_3726(II19373,WX5703,II19371);
  nand NAND2_3727(WX6339,II19372,II19373);
  nand NAND2_3728(II19384,WX5776,WX5705);
  nand NAND2_3729(II19385,WX5776,II19384);
  nand NAND2_3730(II19386,WX5705,II19384);
  nand NAND2_3731(WX6346,II19385,II19386);
  nand NAND2_3732(II19397,WX5777,WX5707);
  nand NAND2_3733(II19398,WX5777,II19397);
  nand NAND2_3734(II19399,WX5707,II19397);
  nand NAND2_3735(WX6353,II19398,II19399);
  nand NAND2_3736(II19410,WX5778,WX5709);
  nand NAND2_3737(II19411,WX5778,II19410);
  nand NAND2_3738(II19412,WX5709,II19410);
  nand NAND2_3739(WX6360,II19411,II19412);
  nand NAND2_3740(II19423,WX5779,WX5711);
  nand NAND2_3741(II19424,WX5779,II19423);
  nand NAND2_3742(II19425,WX5711,II19423);
  nand NAND2_3743(WX6367,II19424,II19425);
  nand NAND2_3744(II19436,WX5780,WX5713);
  nand NAND2_3745(II19437,WX5780,II19436);
  nand NAND2_3746(II19438,WX5713,II19436);
  nand NAND2_3747(WX6374,II19437,II19438);
  nand NAND2_3748(II19449,WX5781,WX5715);
  nand NAND2_3749(II19450,WX5781,II19449);
  nand NAND2_3750(II19451,WX5715,II19449);
  nand NAND2_3751(WX6381,II19450,II19451);
  nand NAND2_3752(II19462,WX5782,WX5717);
  nand NAND2_3753(II19463,WX5782,II19462);
  nand NAND2_3754(II19464,WX5717,II19462);
  nand NAND2_3755(WX6388,II19463,II19464);
  nand NAND2_3756(II19475,WX5783,WX5719);
  nand NAND2_3757(II19476,WX5783,II19475);
  nand NAND2_3758(II19477,WX5719,II19475);
  nand NAND2_3759(WX6395,II19476,II19477);
  nand NAND2_3760(II19490,WX5799,CRC_OUT_5_31);
  nand NAND2_3761(II19491,WX5799,II19490);
  nand NAND2_3762(II19492,CRC_OUT_5_31,II19490);
  nand NAND2_3763(II19489,II19491,II19492);
  nand NAND2_3764(II19497,CRC_OUT_5_15,II19489);
  nand NAND2_3765(II19498,CRC_OUT_5_15,II19497);
  nand NAND2_3766(II19499,II19489,II19497);
  nand NAND2_3767(WX6403,II19498,II19499);
  nand NAND2_3768(II19505,WX5804,CRC_OUT_5_31);
  nand NAND2_3769(II19506,WX5804,II19505);
  nand NAND2_3770(II19507,CRC_OUT_5_31,II19505);
  nand NAND2_3771(II19504,II19506,II19507);
  nand NAND2_3772(II19512,CRC_OUT_5_10,II19504);
  nand NAND2_3773(II19513,CRC_OUT_5_10,II19512);
  nand NAND2_3774(II19514,II19504,II19512);
  nand NAND2_3775(WX6404,II19513,II19514);
  nand NAND2_3776(II19520,WX5811,CRC_OUT_5_31);
  nand NAND2_3777(II19521,WX5811,II19520);
  nand NAND2_3778(II19522,CRC_OUT_5_31,II19520);
  nand NAND2_3779(II19519,II19521,II19522);
  nand NAND2_3780(II19527,CRC_OUT_5_3,II19519);
  nand NAND2_3781(II19528,CRC_OUT_5_3,II19527);
  nand NAND2_3782(II19529,II19519,II19527);
  nand NAND2_3783(WX6405,II19528,II19529);
  nand NAND2_3784(II19534,WX5815,CRC_OUT_5_31);
  nand NAND2_3785(II19535,WX5815,II19534);
  nand NAND2_3786(II19536,CRC_OUT_5_31,II19534);
  nand NAND2_3787(WX6406,II19535,II19536);
  nand NAND2_3788(II19541,WX5784,CRC_OUT_5_30);
  nand NAND2_3789(II19542,WX5784,II19541);
  nand NAND2_3790(II19543,CRC_OUT_5_30,II19541);
  nand NAND2_3791(WX6407,II19542,II19543);
  nand NAND2_3792(II19548,WX5785,CRC_OUT_5_29);
  nand NAND2_3793(II19549,WX5785,II19548);
  nand NAND2_3794(II19550,CRC_OUT_5_29,II19548);
  nand NAND2_3795(WX6408,II19549,II19550);
  nand NAND2_3796(II19555,WX5786,CRC_OUT_5_28);
  nand NAND2_3797(II19556,WX5786,II19555);
  nand NAND2_3798(II19557,CRC_OUT_5_28,II19555);
  nand NAND2_3799(WX6409,II19556,II19557);
  nand NAND2_3800(II19562,WX5787,CRC_OUT_5_27);
  nand NAND2_3801(II19563,WX5787,II19562);
  nand NAND2_3802(II19564,CRC_OUT_5_27,II19562);
  nand NAND2_3803(WX6410,II19563,II19564);
  nand NAND2_3804(II19569,WX5788,CRC_OUT_5_26);
  nand NAND2_3805(II19570,WX5788,II19569);
  nand NAND2_3806(II19571,CRC_OUT_5_26,II19569);
  nand NAND2_3807(WX6411,II19570,II19571);
  nand NAND2_3808(II19576,WX5789,CRC_OUT_5_25);
  nand NAND2_3809(II19577,WX5789,II19576);
  nand NAND2_3810(II19578,CRC_OUT_5_25,II19576);
  nand NAND2_3811(WX6412,II19577,II19578);
  nand NAND2_3812(II19583,WX5790,CRC_OUT_5_24);
  nand NAND2_3813(II19584,WX5790,II19583);
  nand NAND2_3814(II19585,CRC_OUT_5_24,II19583);
  nand NAND2_3815(WX6413,II19584,II19585);
  nand NAND2_3816(II19590,WX5791,CRC_OUT_5_23);
  nand NAND2_3817(II19591,WX5791,II19590);
  nand NAND2_3818(II19592,CRC_OUT_5_23,II19590);
  nand NAND2_3819(WX6414,II19591,II19592);
  nand NAND2_3820(II19597,WX5792,CRC_OUT_5_22);
  nand NAND2_3821(II19598,WX5792,II19597);
  nand NAND2_3822(II19599,CRC_OUT_5_22,II19597);
  nand NAND2_3823(WX6415,II19598,II19599);
  nand NAND2_3824(II19604,WX5793,CRC_OUT_5_21);
  nand NAND2_3825(II19605,WX5793,II19604);
  nand NAND2_3826(II19606,CRC_OUT_5_21,II19604);
  nand NAND2_3827(WX6416,II19605,II19606);
  nand NAND2_3828(II19611,WX5794,CRC_OUT_5_20);
  nand NAND2_3829(II19612,WX5794,II19611);
  nand NAND2_3830(II19613,CRC_OUT_5_20,II19611);
  nand NAND2_3831(WX6417,II19612,II19613);
  nand NAND2_3832(II19618,WX5795,CRC_OUT_5_19);
  nand NAND2_3833(II19619,WX5795,II19618);
  nand NAND2_3834(II19620,CRC_OUT_5_19,II19618);
  nand NAND2_3835(WX6418,II19619,II19620);
  nand NAND2_3836(II19625,WX5796,CRC_OUT_5_18);
  nand NAND2_3837(II19626,WX5796,II19625);
  nand NAND2_3838(II19627,CRC_OUT_5_18,II19625);
  nand NAND2_3839(WX6419,II19626,II19627);
  nand NAND2_3840(II19632,WX5797,CRC_OUT_5_17);
  nand NAND2_3841(II19633,WX5797,II19632);
  nand NAND2_3842(II19634,CRC_OUT_5_17,II19632);
  nand NAND2_3843(WX6420,II19633,II19634);
  nand NAND2_3844(II19639,WX5798,CRC_OUT_5_16);
  nand NAND2_3845(II19640,WX5798,II19639);
  nand NAND2_3846(II19641,CRC_OUT_5_16,II19639);
  nand NAND2_3847(WX6421,II19640,II19641);
  nand NAND2_3848(II19646,WX5800,CRC_OUT_5_14);
  nand NAND2_3849(II19647,WX5800,II19646);
  nand NAND2_3850(II19648,CRC_OUT_5_14,II19646);
  nand NAND2_3851(WX6422,II19647,II19648);
  nand NAND2_3852(II19653,WX5801,CRC_OUT_5_13);
  nand NAND2_3853(II19654,WX5801,II19653);
  nand NAND2_3854(II19655,CRC_OUT_5_13,II19653);
  nand NAND2_3855(WX6423,II19654,II19655);
  nand NAND2_3856(II19660,WX5802,CRC_OUT_5_12);
  nand NAND2_3857(II19661,WX5802,II19660);
  nand NAND2_3858(II19662,CRC_OUT_5_12,II19660);
  nand NAND2_3859(WX6424,II19661,II19662);
  nand NAND2_3860(II19667,WX5803,CRC_OUT_5_11);
  nand NAND2_3861(II19668,WX5803,II19667);
  nand NAND2_3862(II19669,CRC_OUT_5_11,II19667);
  nand NAND2_3863(WX6425,II19668,II19669);
  nand NAND2_3864(II19674,WX5805,CRC_OUT_5_9);
  nand NAND2_3865(II19675,WX5805,II19674);
  nand NAND2_3866(II19676,CRC_OUT_5_9,II19674);
  nand NAND2_3867(WX6426,II19675,II19676);
  nand NAND2_3868(II19681,WX5806,CRC_OUT_5_8);
  nand NAND2_3869(II19682,WX5806,II19681);
  nand NAND2_3870(II19683,CRC_OUT_5_8,II19681);
  nand NAND2_3871(WX6427,II19682,II19683);
  nand NAND2_3872(II19688,WX5807,CRC_OUT_5_7);
  nand NAND2_3873(II19689,WX5807,II19688);
  nand NAND2_3874(II19690,CRC_OUT_5_7,II19688);
  nand NAND2_3875(WX6428,II19689,II19690);
  nand NAND2_3876(II19695,WX5808,CRC_OUT_5_6);
  nand NAND2_3877(II19696,WX5808,II19695);
  nand NAND2_3878(II19697,CRC_OUT_5_6,II19695);
  nand NAND2_3879(WX6429,II19696,II19697);
  nand NAND2_3880(II19702,WX5809,CRC_OUT_5_5);
  nand NAND2_3881(II19703,WX5809,II19702);
  nand NAND2_3882(II19704,CRC_OUT_5_5,II19702);
  nand NAND2_3883(WX6430,II19703,II19704);
  nand NAND2_3884(II19709,WX5810,CRC_OUT_5_4);
  nand NAND2_3885(II19710,WX5810,II19709);
  nand NAND2_3886(II19711,CRC_OUT_5_4,II19709);
  nand NAND2_3887(WX6431,II19710,II19711);
  nand NAND2_3888(II19716,WX5812,CRC_OUT_5_2);
  nand NAND2_3889(II19717,WX5812,II19716);
  nand NAND2_3890(II19718,CRC_OUT_5_2,II19716);
  nand NAND2_3891(WX6432,II19717,II19718);
  nand NAND2_3892(II19723,WX5813,CRC_OUT_5_1);
  nand NAND2_3893(II19724,WX5813,II19723);
  nand NAND2_3894(II19725,CRC_OUT_5_1,II19723);
  nand NAND2_3895(WX6433,II19724,II19725);
  nand NAND2_3896(II19730,WX5814,CRC_OUT_5_0);
  nand NAND2_3897(II19731,WX5814,II19730);
  nand NAND2_3898(II19732,CRC_OUT_5_0,II19730);
  nand NAND2_3899(WX6434,II19731,II19732);
  nand NAND2_3900(II22013,WX7466,WX7110);
  nand NAND2_3901(II22014,WX7466,II22013);
  nand NAND2_3902(II22015,WX7110,II22013);
  nand NAND2_3903(II22012,II22014,II22015);
  nand NAND2_3904(II22020,WX7174,II22012);
  nand NAND2_3905(II22021,WX7174,II22020);
  nand NAND2_3906(II22022,II22012,II22020);
  nand NAND2_3907(II22011,II22021,II22022);
  nand NAND2_3908(II22028,WX7238,WX7302);
  nand NAND2_3909(II22029,WX7238,II22028);
  nand NAND2_3910(II22030,WX7302,II22028);
  nand NAND2_3911(II22027,II22029,II22030);
  nand NAND2_3912(II22035,II22011,II22027);
  nand NAND2_3913(II22036,II22011,II22035);
  nand NAND2_3914(II22037,II22027,II22035);
  nand NAND2_3915(WX7365,II22036,II22037);
  nand NAND2_3916(II22044,WX7466,WX7112);
  nand NAND2_3917(II22045,WX7466,II22044);
  nand NAND2_3918(II22046,WX7112,II22044);
  nand NAND2_3919(II22043,II22045,II22046);
  nand NAND2_3920(II22051,WX7176,II22043);
  nand NAND2_3921(II22052,WX7176,II22051);
  nand NAND2_3922(II22053,II22043,II22051);
  nand NAND2_3923(II22042,II22052,II22053);
  nand NAND2_3924(II22059,WX7240,WX7304);
  nand NAND2_3925(II22060,WX7240,II22059);
  nand NAND2_3926(II22061,WX7304,II22059);
  nand NAND2_3927(II22058,II22060,II22061);
  nand NAND2_3928(II22066,II22042,II22058);
  nand NAND2_3929(II22067,II22042,II22066);
  nand NAND2_3930(II22068,II22058,II22066);
  nand NAND2_3931(WX7366,II22067,II22068);
  nand NAND2_3932(II22075,WX7466,WX7114);
  nand NAND2_3933(II22076,WX7466,II22075);
  nand NAND2_3934(II22077,WX7114,II22075);
  nand NAND2_3935(II22074,II22076,II22077);
  nand NAND2_3936(II22082,WX7178,II22074);
  nand NAND2_3937(II22083,WX7178,II22082);
  nand NAND2_3938(II22084,II22074,II22082);
  nand NAND2_3939(II22073,II22083,II22084);
  nand NAND2_3940(II22090,WX7242,WX7306);
  nand NAND2_3941(II22091,WX7242,II22090);
  nand NAND2_3942(II22092,WX7306,II22090);
  nand NAND2_3943(II22089,II22091,II22092);
  nand NAND2_3944(II22097,II22073,II22089);
  nand NAND2_3945(II22098,II22073,II22097);
  nand NAND2_3946(II22099,II22089,II22097);
  nand NAND2_3947(WX7367,II22098,II22099);
  nand NAND2_3948(II22106,WX7466,WX7116);
  nand NAND2_3949(II22107,WX7466,II22106);
  nand NAND2_3950(II22108,WX7116,II22106);
  nand NAND2_3951(II22105,II22107,II22108);
  nand NAND2_3952(II22113,WX7180,II22105);
  nand NAND2_3953(II22114,WX7180,II22113);
  nand NAND2_3954(II22115,II22105,II22113);
  nand NAND2_3955(II22104,II22114,II22115);
  nand NAND2_3956(II22121,WX7244,WX7308);
  nand NAND2_3957(II22122,WX7244,II22121);
  nand NAND2_3958(II22123,WX7308,II22121);
  nand NAND2_3959(II22120,II22122,II22123);
  nand NAND2_3960(II22128,II22104,II22120);
  nand NAND2_3961(II22129,II22104,II22128);
  nand NAND2_3962(II22130,II22120,II22128);
  nand NAND2_3963(WX7368,II22129,II22130);
  nand NAND2_3964(II22137,WX7466,WX7118);
  nand NAND2_3965(II22138,WX7466,II22137);
  nand NAND2_3966(II22139,WX7118,II22137);
  nand NAND2_3967(II22136,II22138,II22139);
  nand NAND2_3968(II22144,WX7182,II22136);
  nand NAND2_3969(II22145,WX7182,II22144);
  nand NAND2_3970(II22146,II22136,II22144);
  nand NAND2_3971(II22135,II22145,II22146);
  nand NAND2_3972(II22152,WX7246,WX7310);
  nand NAND2_3973(II22153,WX7246,II22152);
  nand NAND2_3974(II22154,WX7310,II22152);
  nand NAND2_3975(II22151,II22153,II22154);
  nand NAND2_3976(II22159,II22135,II22151);
  nand NAND2_3977(II22160,II22135,II22159);
  nand NAND2_3978(II22161,II22151,II22159);
  nand NAND2_3979(WX7369,II22160,II22161);
  nand NAND2_3980(II22168,WX7466,WX7120);
  nand NAND2_3981(II22169,WX7466,II22168);
  nand NAND2_3982(II22170,WX7120,II22168);
  nand NAND2_3983(II22167,II22169,II22170);
  nand NAND2_3984(II22175,WX7184,II22167);
  nand NAND2_3985(II22176,WX7184,II22175);
  nand NAND2_3986(II22177,II22167,II22175);
  nand NAND2_3987(II22166,II22176,II22177);
  nand NAND2_3988(II22183,WX7248,WX7312);
  nand NAND2_3989(II22184,WX7248,II22183);
  nand NAND2_3990(II22185,WX7312,II22183);
  nand NAND2_3991(II22182,II22184,II22185);
  nand NAND2_3992(II22190,II22166,II22182);
  nand NAND2_3993(II22191,II22166,II22190);
  nand NAND2_3994(II22192,II22182,II22190);
  nand NAND2_3995(WX7370,II22191,II22192);
  nand NAND2_3996(II22199,WX7466,WX7122);
  nand NAND2_3997(II22200,WX7466,II22199);
  nand NAND2_3998(II22201,WX7122,II22199);
  nand NAND2_3999(II22198,II22200,II22201);
  nand NAND2_4000(II22206,WX7186,II22198);
  nand NAND2_4001(II22207,WX7186,II22206);
  nand NAND2_4002(II22208,II22198,II22206);
  nand NAND2_4003(II22197,II22207,II22208);
  nand NAND2_4004(II22214,WX7250,WX7314);
  nand NAND2_4005(II22215,WX7250,II22214);
  nand NAND2_4006(II22216,WX7314,II22214);
  nand NAND2_4007(II22213,II22215,II22216);
  nand NAND2_4008(II22221,II22197,II22213);
  nand NAND2_4009(II22222,II22197,II22221);
  nand NAND2_4010(II22223,II22213,II22221);
  nand NAND2_4011(WX7371,II22222,II22223);
  nand NAND2_4012(II22230,WX7466,WX7124);
  nand NAND2_4013(II22231,WX7466,II22230);
  nand NAND2_4014(II22232,WX7124,II22230);
  nand NAND2_4015(II22229,II22231,II22232);
  nand NAND2_4016(II22237,WX7188,II22229);
  nand NAND2_4017(II22238,WX7188,II22237);
  nand NAND2_4018(II22239,II22229,II22237);
  nand NAND2_4019(II22228,II22238,II22239);
  nand NAND2_4020(II22245,WX7252,WX7316);
  nand NAND2_4021(II22246,WX7252,II22245);
  nand NAND2_4022(II22247,WX7316,II22245);
  nand NAND2_4023(II22244,II22246,II22247);
  nand NAND2_4024(II22252,II22228,II22244);
  nand NAND2_4025(II22253,II22228,II22252);
  nand NAND2_4026(II22254,II22244,II22252);
  nand NAND2_4027(WX7372,II22253,II22254);
  nand NAND2_4028(II22261,WX7466,WX7126);
  nand NAND2_4029(II22262,WX7466,II22261);
  nand NAND2_4030(II22263,WX7126,II22261);
  nand NAND2_4031(II22260,II22262,II22263);
  nand NAND2_4032(II22268,WX7190,II22260);
  nand NAND2_4033(II22269,WX7190,II22268);
  nand NAND2_4034(II22270,II22260,II22268);
  nand NAND2_4035(II22259,II22269,II22270);
  nand NAND2_4036(II22276,WX7254,WX7318);
  nand NAND2_4037(II22277,WX7254,II22276);
  nand NAND2_4038(II22278,WX7318,II22276);
  nand NAND2_4039(II22275,II22277,II22278);
  nand NAND2_4040(II22283,II22259,II22275);
  nand NAND2_4041(II22284,II22259,II22283);
  nand NAND2_4042(II22285,II22275,II22283);
  nand NAND2_4043(WX7373,II22284,II22285);
  nand NAND2_4044(II22292,WX7466,WX7128);
  nand NAND2_4045(II22293,WX7466,II22292);
  nand NAND2_4046(II22294,WX7128,II22292);
  nand NAND2_4047(II22291,II22293,II22294);
  nand NAND2_4048(II22299,WX7192,II22291);
  nand NAND2_4049(II22300,WX7192,II22299);
  nand NAND2_4050(II22301,II22291,II22299);
  nand NAND2_4051(II22290,II22300,II22301);
  nand NAND2_4052(II22307,WX7256,WX7320);
  nand NAND2_4053(II22308,WX7256,II22307);
  nand NAND2_4054(II22309,WX7320,II22307);
  nand NAND2_4055(II22306,II22308,II22309);
  nand NAND2_4056(II22314,II22290,II22306);
  nand NAND2_4057(II22315,II22290,II22314);
  nand NAND2_4058(II22316,II22306,II22314);
  nand NAND2_4059(WX7374,II22315,II22316);
  nand NAND2_4060(II22323,WX7466,WX7130);
  nand NAND2_4061(II22324,WX7466,II22323);
  nand NAND2_4062(II22325,WX7130,II22323);
  nand NAND2_4063(II22322,II22324,II22325);
  nand NAND2_4064(II22330,WX7194,II22322);
  nand NAND2_4065(II22331,WX7194,II22330);
  nand NAND2_4066(II22332,II22322,II22330);
  nand NAND2_4067(II22321,II22331,II22332);
  nand NAND2_4068(II22338,WX7258,WX7322);
  nand NAND2_4069(II22339,WX7258,II22338);
  nand NAND2_4070(II22340,WX7322,II22338);
  nand NAND2_4071(II22337,II22339,II22340);
  nand NAND2_4072(II22345,II22321,II22337);
  nand NAND2_4073(II22346,II22321,II22345);
  nand NAND2_4074(II22347,II22337,II22345);
  nand NAND2_4075(WX7375,II22346,II22347);
  nand NAND2_4076(II22354,WX7466,WX7132);
  nand NAND2_4077(II22355,WX7466,II22354);
  nand NAND2_4078(II22356,WX7132,II22354);
  nand NAND2_4079(II22353,II22355,II22356);
  nand NAND2_4080(II22361,WX7196,II22353);
  nand NAND2_4081(II22362,WX7196,II22361);
  nand NAND2_4082(II22363,II22353,II22361);
  nand NAND2_4083(II22352,II22362,II22363);
  nand NAND2_4084(II22369,WX7260,WX7324);
  nand NAND2_4085(II22370,WX7260,II22369);
  nand NAND2_4086(II22371,WX7324,II22369);
  nand NAND2_4087(II22368,II22370,II22371);
  nand NAND2_4088(II22376,II22352,II22368);
  nand NAND2_4089(II22377,II22352,II22376);
  nand NAND2_4090(II22378,II22368,II22376);
  nand NAND2_4091(WX7376,II22377,II22378);
  nand NAND2_4092(II22385,WX7466,WX7134);
  nand NAND2_4093(II22386,WX7466,II22385);
  nand NAND2_4094(II22387,WX7134,II22385);
  nand NAND2_4095(II22384,II22386,II22387);
  nand NAND2_4096(II22392,WX7198,II22384);
  nand NAND2_4097(II22393,WX7198,II22392);
  nand NAND2_4098(II22394,II22384,II22392);
  nand NAND2_4099(II22383,II22393,II22394);
  nand NAND2_4100(II22400,WX7262,WX7326);
  nand NAND2_4101(II22401,WX7262,II22400);
  nand NAND2_4102(II22402,WX7326,II22400);
  nand NAND2_4103(II22399,II22401,II22402);
  nand NAND2_4104(II22407,II22383,II22399);
  nand NAND2_4105(II22408,II22383,II22407);
  nand NAND2_4106(II22409,II22399,II22407);
  nand NAND2_4107(WX7377,II22408,II22409);
  nand NAND2_4108(II22416,WX7466,WX7136);
  nand NAND2_4109(II22417,WX7466,II22416);
  nand NAND2_4110(II22418,WX7136,II22416);
  nand NAND2_4111(II22415,II22417,II22418);
  nand NAND2_4112(II22423,WX7200,II22415);
  nand NAND2_4113(II22424,WX7200,II22423);
  nand NAND2_4114(II22425,II22415,II22423);
  nand NAND2_4115(II22414,II22424,II22425);
  nand NAND2_4116(II22431,WX7264,WX7328);
  nand NAND2_4117(II22432,WX7264,II22431);
  nand NAND2_4118(II22433,WX7328,II22431);
  nand NAND2_4119(II22430,II22432,II22433);
  nand NAND2_4120(II22438,II22414,II22430);
  nand NAND2_4121(II22439,II22414,II22438);
  nand NAND2_4122(II22440,II22430,II22438);
  nand NAND2_4123(WX7378,II22439,II22440);
  nand NAND2_4124(II22447,WX7466,WX7138);
  nand NAND2_4125(II22448,WX7466,II22447);
  nand NAND2_4126(II22449,WX7138,II22447);
  nand NAND2_4127(II22446,II22448,II22449);
  nand NAND2_4128(II22454,WX7202,II22446);
  nand NAND2_4129(II22455,WX7202,II22454);
  nand NAND2_4130(II22456,II22446,II22454);
  nand NAND2_4131(II22445,II22455,II22456);
  nand NAND2_4132(II22462,WX7266,WX7330);
  nand NAND2_4133(II22463,WX7266,II22462);
  nand NAND2_4134(II22464,WX7330,II22462);
  nand NAND2_4135(II22461,II22463,II22464);
  nand NAND2_4136(II22469,II22445,II22461);
  nand NAND2_4137(II22470,II22445,II22469);
  nand NAND2_4138(II22471,II22461,II22469);
  nand NAND2_4139(WX7379,II22470,II22471);
  nand NAND2_4140(II22478,WX7466,WX7140);
  nand NAND2_4141(II22479,WX7466,II22478);
  nand NAND2_4142(II22480,WX7140,II22478);
  nand NAND2_4143(II22477,II22479,II22480);
  nand NAND2_4144(II22485,WX7204,II22477);
  nand NAND2_4145(II22486,WX7204,II22485);
  nand NAND2_4146(II22487,II22477,II22485);
  nand NAND2_4147(II22476,II22486,II22487);
  nand NAND2_4148(II22493,WX7268,WX7332);
  nand NAND2_4149(II22494,WX7268,II22493);
  nand NAND2_4150(II22495,WX7332,II22493);
  nand NAND2_4151(II22492,II22494,II22495);
  nand NAND2_4152(II22500,II22476,II22492);
  nand NAND2_4153(II22501,II22476,II22500);
  nand NAND2_4154(II22502,II22492,II22500);
  nand NAND2_4155(WX7380,II22501,II22502);
  nand NAND2_4156(II22509,WX7467,WX7142);
  nand NAND2_4157(II22510,WX7467,II22509);
  nand NAND2_4158(II22511,WX7142,II22509);
  nand NAND2_4159(II22508,II22510,II22511);
  nand NAND2_4160(II22516,WX7206,II22508);
  nand NAND2_4161(II22517,WX7206,II22516);
  nand NAND2_4162(II22518,II22508,II22516);
  nand NAND2_4163(II22507,II22517,II22518);
  nand NAND2_4164(II22524,WX7270,WX7334);
  nand NAND2_4165(II22525,WX7270,II22524);
  nand NAND2_4166(II22526,WX7334,II22524);
  nand NAND2_4167(II22523,II22525,II22526);
  nand NAND2_4168(II22531,II22507,II22523);
  nand NAND2_4169(II22532,II22507,II22531);
  nand NAND2_4170(II22533,II22523,II22531);
  nand NAND2_4171(WX7381,II22532,II22533);
  nand NAND2_4172(II22540,WX7467,WX7144);
  nand NAND2_4173(II22541,WX7467,II22540);
  nand NAND2_4174(II22542,WX7144,II22540);
  nand NAND2_4175(II22539,II22541,II22542);
  nand NAND2_4176(II22547,WX7208,II22539);
  nand NAND2_4177(II22548,WX7208,II22547);
  nand NAND2_4178(II22549,II22539,II22547);
  nand NAND2_4179(II22538,II22548,II22549);
  nand NAND2_4180(II22555,WX7272,WX7336);
  nand NAND2_4181(II22556,WX7272,II22555);
  nand NAND2_4182(II22557,WX7336,II22555);
  nand NAND2_4183(II22554,II22556,II22557);
  nand NAND2_4184(II22562,II22538,II22554);
  nand NAND2_4185(II22563,II22538,II22562);
  nand NAND2_4186(II22564,II22554,II22562);
  nand NAND2_4187(WX7382,II22563,II22564);
  nand NAND2_4188(II22571,WX7467,WX7146);
  nand NAND2_4189(II22572,WX7467,II22571);
  nand NAND2_4190(II22573,WX7146,II22571);
  nand NAND2_4191(II22570,II22572,II22573);
  nand NAND2_4192(II22578,WX7210,II22570);
  nand NAND2_4193(II22579,WX7210,II22578);
  nand NAND2_4194(II22580,II22570,II22578);
  nand NAND2_4195(II22569,II22579,II22580);
  nand NAND2_4196(II22586,WX7274,WX7338);
  nand NAND2_4197(II22587,WX7274,II22586);
  nand NAND2_4198(II22588,WX7338,II22586);
  nand NAND2_4199(II22585,II22587,II22588);
  nand NAND2_4200(II22593,II22569,II22585);
  nand NAND2_4201(II22594,II22569,II22593);
  nand NAND2_4202(II22595,II22585,II22593);
  nand NAND2_4203(WX7383,II22594,II22595);
  nand NAND2_4204(II22602,WX7467,WX7148);
  nand NAND2_4205(II22603,WX7467,II22602);
  nand NAND2_4206(II22604,WX7148,II22602);
  nand NAND2_4207(II22601,II22603,II22604);
  nand NAND2_4208(II22609,WX7212,II22601);
  nand NAND2_4209(II22610,WX7212,II22609);
  nand NAND2_4210(II22611,II22601,II22609);
  nand NAND2_4211(II22600,II22610,II22611);
  nand NAND2_4212(II22617,WX7276,WX7340);
  nand NAND2_4213(II22618,WX7276,II22617);
  nand NAND2_4214(II22619,WX7340,II22617);
  nand NAND2_4215(II22616,II22618,II22619);
  nand NAND2_4216(II22624,II22600,II22616);
  nand NAND2_4217(II22625,II22600,II22624);
  nand NAND2_4218(II22626,II22616,II22624);
  nand NAND2_4219(WX7384,II22625,II22626);
  nand NAND2_4220(II22633,WX7467,WX7150);
  nand NAND2_4221(II22634,WX7467,II22633);
  nand NAND2_4222(II22635,WX7150,II22633);
  nand NAND2_4223(II22632,II22634,II22635);
  nand NAND2_4224(II22640,WX7214,II22632);
  nand NAND2_4225(II22641,WX7214,II22640);
  nand NAND2_4226(II22642,II22632,II22640);
  nand NAND2_4227(II22631,II22641,II22642);
  nand NAND2_4228(II22648,WX7278,WX7342);
  nand NAND2_4229(II22649,WX7278,II22648);
  nand NAND2_4230(II22650,WX7342,II22648);
  nand NAND2_4231(II22647,II22649,II22650);
  nand NAND2_4232(II22655,II22631,II22647);
  nand NAND2_4233(II22656,II22631,II22655);
  nand NAND2_4234(II22657,II22647,II22655);
  nand NAND2_4235(WX7385,II22656,II22657);
  nand NAND2_4236(II22664,WX7467,WX7152);
  nand NAND2_4237(II22665,WX7467,II22664);
  nand NAND2_4238(II22666,WX7152,II22664);
  nand NAND2_4239(II22663,II22665,II22666);
  nand NAND2_4240(II22671,WX7216,II22663);
  nand NAND2_4241(II22672,WX7216,II22671);
  nand NAND2_4242(II22673,II22663,II22671);
  nand NAND2_4243(II22662,II22672,II22673);
  nand NAND2_4244(II22679,WX7280,WX7344);
  nand NAND2_4245(II22680,WX7280,II22679);
  nand NAND2_4246(II22681,WX7344,II22679);
  nand NAND2_4247(II22678,II22680,II22681);
  nand NAND2_4248(II22686,II22662,II22678);
  nand NAND2_4249(II22687,II22662,II22686);
  nand NAND2_4250(II22688,II22678,II22686);
  nand NAND2_4251(WX7386,II22687,II22688);
  nand NAND2_4252(II22695,WX7467,WX7154);
  nand NAND2_4253(II22696,WX7467,II22695);
  nand NAND2_4254(II22697,WX7154,II22695);
  nand NAND2_4255(II22694,II22696,II22697);
  nand NAND2_4256(II22702,WX7218,II22694);
  nand NAND2_4257(II22703,WX7218,II22702);
  nand NAND2_4258(II22704,II22694,II22702);
  nand NAND2_4259(II22693,II22703,II22704);
  nand NAND2_4260(II22710,WX7282,WX7346);
  nand NAND2_4261(II22711,WX7282,II22710);
  nand NAND2_4262(II22712,WX7346,II22710);
  nand NAND2_4263(II22709,II22711,II22712);
  nand NAND2_4264(II22717,II22693,II22709);
  nand NAND2_4265(II22718,II22693,II22717);
  nand NAND2_4266(II22719,II22709,II22717);
  nand NAND2_4267(WX7387,II22718,II22719);
  nand NAND2_4268(II22726,WX7467,WX7156);
  nand NAND2_4269(II22727,WX7467,II22726);
  nand NAND2_4270(II22728,WX7156,II22726);
  nand NAND2_4271(II22725,II22727,II22728);
  nand NAND2_4272(II22733,WX7220,II22725);
  nand NAND2_4273(II22734,WX7220,II22733);
  nand NAND2_4274(II22735,II22725,II22733);
  nand NAND2_4275(II22724,II22734,II22735);
  nand NAND2_4276(II22741,WX7284,WX7348);
  nand NAND2_4277(II22742,WX7284,II22741);
  nand NAND2_4278(II22743,WX7348,II22741);
  nand NAND2_4279(II22740,II22742,II22743);
  nand NAND2_4280(II22748,II22724,II22740);
  nand NAND2_4281(II22749,II22724,II22748);
  nand NAND2_4282(II22750,II22740,II22748);
  nand NAND2_4283(WX7388,II22749,II22750);
  nand NAND2_4284(II22757,WX7467,WX7158);
  nand NAND2_4285(II22758,WX7467,II22757);
  nand NAND2_4286(II22759,WX7158,II22757);
  nand NAND2_4287(II22756,II22758,II22759);
  nand NAND2_4288(II22764,WX7222,II22756);
  nand NAND2_4289(II22765,WX7222,II22764);
  nand NAND2_4290(II22766,II22756,II22764);
  nand NAND2_4291(II22755,II22765,II22766);
  nand NAND2_4292(II22772,WX7286,WX7350);
  nand NAND2_4293(II22773,WX7286,II22772);
  nand NAND2_4294(II22774,WX7350,II22772);
  nand NAND2_4295(II22771,II22773,II22774);
  nand NAND2_4296(II22779,II22755,II22771);
  nand NAND2_4297(II22780,II22755,II22779);
  nand NAND2_4298(II22781,II22771,II22779);
  nand NAND2_4299(WX7389,II22780,II22781);
  nand NAND2_4300(II22788,WX7467,WX7160);
  nand NAND2_4301(II22789,WX7467,II22788);
  nand NAND2_4302(II22790,WX7160,II22788);
  nand NAND2_4303(II22787,II22789,II22790);
  nand NAND2_4304(II22795,WX7224,II22787);
  nand NAND2_4305(II22796,WX7224,II22795);
  nand NAND2_4306(II22797,II22787,II22795);
  nand NAND2_4307(II22786,II22796,II22797);
  nand NAND2_4308(II22803,WX7288,WX7352);
  nand NAND2_4309(II22804,WX7288,II22803);
  nand NAND2_4310(II22805,WX7352,II22803);
  nand NAND2_4311(II22802,II22804,II22805);
  nand NAND2_4312(II22810,II22786,II22802);
  nand NAND2_4313(II22811,II22786,II22810);
  nand NAND2_4314(II22812,II22802,II22810);
  nand NAND2_4315(WX7390,II22811,II22812);
  nand NAND2_4316(II22819,WX7467,WX7162);
  nand NAND2_4317(II22820,WX7467,II22819);
  nand NAND2_4318(II22821,WX7162,II22819);
  nand NAND2_4319(II22818,II22820,II22821);
  nand NAND2_4320(II22826,WX7226,II22818);
  nand NAND2_4321(II22827,WX7226,II22826);
  nand NAND2_4322(II22828,II22818,II22826);
  nand NAND2_4323(II22817,II22827,II22828);
  nand NAND2_4324(II22834,WX7290,WX7354);
  nand NAND2_4325(II22835,WX7290,II22834);
  nand NAND2_4326(II22836,WX7354,II22834);
  nand NAND2_4327(II22833,II22835,II22836);
  nand NAND2_4328(II22841,II22817,II22833);
  nand NAND2_4329(II22842,II22817,II22841);
  nand NAND2_4330(II22843,II22833,II22841);
  nand NAND2_4331(WX7391,II22842,II22843);
  nand NAND2_4332(II22850,WX7467,WX7164);
  nand NAND2_4333(II22851,WX7467,II22850);
  nand NAND2_4334(II22852,WX7164,II22850);
  nand NAND2_4335(II22849,II22851,II22852);
  nand NAND2_4336(II22857,WX7228,II22849);
  nand NAND2_4337(II22858,WX7228,II22857);
  nand NAND2_4338(II22859,II22849,II22857);
  nand NAND2_4339(II22848,II22858,II22859);
  nand NAND2_4340(II22865,WX7292,WX7356);
  nand NAND2_4341(II22866,WX7292,II22865);
  nand NAND2_4342(II22867,WX7356,II22865);
  nand NAND2_4343(II22864,II22866,II22867);
  nand NAND2_4344(II22872,II22848,II22864);
  nand NAND2_4345(II22873,II22848,II22872);
  nand NAND2_4346(II22874,II22864,II22872);
  nand NAND2_4347(WX7392,II22873,II22874);
  nand NAND2_4348(II22881,WX7467,WX7166);
  nand NAND2_4349(II22882,WX7467,II22881);
  nand NAND2_4350(II22883,WX7166,II22881);
  nand NAND2_4351(II22880,II22882,II22883);
  nand NAND2_4352(II22888,WX7230,II22880);
  nand NAND2_4353(II22889,WX7230,II22888);
  nand NAND2_4354(II22890,II22880,II22888);
  nand NAND2_4355(II22879,II22889,II22890);
  nand NAND2_4356(II22896,WX7294,WX7358);
  nand NAND2_4357(II22897,WX7294,II22896);
  nand NAND2_4358(II22898,WX7358,II22896);
  nand NAND2_4359(II22895,II22897,II22898);
  nand NAND2_4360(II22903,II22879,II22895);
  nand NAND2_4361(II22904,II22879,II22903);
  nand NAND2_4362(II22905,II22895,II22903);
  nand NAND2_4363(WX7393,II22904,II22905);
  nand NAND2_4364(II22912,WX7467,WX7168);
  nand NAND2_4365(II22913,WX7467,II22912);
  nand NAND2_4366(II22914,WX7168,II22912);
  nand NAND2_4367(II22911,II22913,II22914);
  nand NAND2_4368(II22919,WX7232,II22911);
  nand NAND2_4369(II22920,WX7232,II22919);
  nand NAND2_4370(II22921,II22911,II22919);
  nand NAND2_4371(II22910,II22920,II22921);
  nand NAND2_4372(II22927,WX7296,WX7360);
  nand NAND2_4373(II22928,WX7296,II22927);
  nand NAND2_4374(II22929,WX7360,II22927);
  nand NAND2_4375(II22926,II22928,II22929);
  nand NAND2_4376(II22934,II22910,II22926);
  nand NAND2_4377(II22935,II22910,II22934);
  nand NAND2_4378(II22936,II22926,II22934);
  nand NAND2_4379(WX7394,II22935,II22936);
  nand NAND2_4380(II22943,WX7467,WX7170);
  nand NAND2_4381(II22944,WX7467,II22943);
  nand NAND2_4382(II22945,WX7170,II22943);
  nand NAND2_4383(II22942,II22944,II22945);
  nand NAND2_4384(II22950,WX7234,II22942);
  nand NAND2_4385(II22951,WX7234,II22950);
  nand NAND2_4386(II22952,II22942,II22950);
  nand NAND2_4387(II22941,II22951,II22952);
  nand NAND2_4388(II22958,WX7298,WX7362);
  nand NAND2_4389(II22959,WX7298,II22958);
  nand NAND2_4390(II22960,WX7362,II22958);
  nand NAND2_4391(II22957,II22959,II22960);
  nand NAND2_4392(II22965,II22941,II22957);
  nand NAND2_4393(II22966,II22941,II22965);
  nand NAND2_4394(II22967,II22957,II22965);
  nand NAND2_4395(WX7395,II22966,II22967);
  nand NAND2_4396(II22974,WX7467,WX7172);
  nand NAND2_4397(II22975,WX7467,II22974);
  nand NAND2_4398(II22976,WX7172,II22974);
  nand NAND2_4399(II22973,II22975,II22976);
  nand NAND2_4400(II22981,WX7236,II22973);
  nand NAND2_4401(II22982,WX7236,II22981);
  nand NAND2_4402(II22983,II22973,II22981);
  nand NAND2_4403(II22972,II22982,II22983);
  nand NAND2_4404(II22989,WX7300,WX7364);
  nand NAND2_4405(II22990,WX7300,II22989);
  nand NAND2_4406(II22991,WX7364,II22989);
  nand NAND2_4407(II22988,II22990,II22991);
  nand NAND2_4408(II22996,II22972,II22988);
  nand NAND2_4409(II22997,II22972,II22996);
  nand NAND2_4410(II22998,II22988,II22996);
  nand NAND2_4411(WX7396,II22997,II22998);
  nand NAND2_4412(II23077,WX7045,WX6950);
  nand NAND2_4413(II23078,WX7045,II23077);
  nand NAND2_4414(II23079,WX6950,II23077);
  nand NAND2_4415(WX7471,II23078,II23079);
  nand NAND2_4416(II23090,WX7046,WX6952);
  nand NAND2_4417(II23091,WX7046,II23090);
  nand NAND2_4418(II23092,WX6952,II23090);
  nand NAND2_4419(WX7478,II23091,II23092);
  nand NAND2_4420(II23103,WX7047,WX6954);
  nand NAND2_4421(II23104,WX7047,II23103);
  nand NAND2_4422(II23105,WX6954,II23103);
  nand NAND2_4423(WX7485,II23104,II23105);
  nand NAND2_4424(II23116,WX7048,WX6956);
  nand NAND2_4425(II23117,WX7048,II23116);
  nand NAND2_4426(II23118,WX6956,II23116);
  nand NAND2_4427(WX7492,II23117,II23118);
  nand NAND2_4428(II23129,WX7049,WX6958);
  nand NAND2_4429(II23130,WX7049,II23129);
  nand NAND2_4430(II23131,WX6958,II23129);
  nand NAND2_4431(WX7499,II23130,II23131);
  nand NAND2_4432(II23142,WX7050,WX6960);
  nand NAND2_4433(II23143,WX7050,II23142);
  nand NAND2_4434(II23144,WX6960,II23142);
  nand NAND2_4435(WX7506,II23143,II23144);
  nand NAND2_4436(II23155,WX7051,WX6962);
  nand NAND2_4437(II23156,WX7051,II23155);
  nand NAND2_4438(II23157,WX6962,II23155);
  nand NAND2_4439(WX7513,II23156,II23157);
  nand NAND2_4440(II23168,WX7052,WX6964);
  nand NAND2_4441(II23169,WX7052,II23168);
  nand NAND2_4442(II23170,WX6964,II23168);
  nand NAND2_4443(WX7520,II23169,II23170);
  nand NAND2_4444(II23181,WX7053,WX6966);
  nand NAND2_4445(II23182,WX7053,II23181);
  nand NAND2_4446(II23183,WX6966,II23181);
  nand NAND2_4447(WX7527,II23182,II23183);
  nand NAND2_4448(II23194,WX7054,WX6968);
  nand NAND2_4449(II23195,WX7054,II23194);
  nand NAND2_4450(II23196,WX6968,II23194);
  nand NAND2_4451(WX7534,II23195,II23196);
  nand NAND2_4452(II23207,WX7055,WX6970);
  nand NAND2_4453(II23208,WX7055,II23207);
  nand NAND2_4454(II23209,WX6970,II23207);
  nand NAND2_4455(WX7541,II23208,II23209);
  nand NAND2_4456(II23220,WX7056,WX6972);
  nand NAND2_4457(II23221,WX7056,II23220);
  nand NAND2_4458(II23222,WX6972,II23220);
  nand NAND2_4459(WX7548,II23221,II23222);
  nand NAND2_4460(II23233,WX7057,WX6974);
  nand NAND2_4461(II23234,WX7057,II23233);
  nand NAND2_4462(II23235,WX6974,II23233);
  nand NAND2_4463(WX7555,II23234,II23235);
  nand NAND2_4464(II23246,WX7058,WX6976);
  nand NAND2_4465(II23247,WX7058,II23246);
  nand NAND2_4466(II23248,WX6976,II23246);
  nand NAND2_4467(WX7562,II23247,II23248);
  nand NAND2_4468(II23259,WX7059,WX6978);
  nand NAND2_4469(II23260,WX7059,II23259);
  nand NAND2_4470(II23261,WX6978,II23259);
  nand NAND2_4471(WX7569,II23260,II23261);
  nand NAND2_4472(II23272,WX7060,WX6980);
  nand NAND2_4473(II23273,WX7060,II23272);
  nand NAND2_4474(II23274,WX6980,II23272);
  nand NAND2_4475(WX7576,II23273,II23274);
  nand NAND2_4476(II23285,WX7061,WX6982);
  nand NAND2_4477(II23286,WX7061,II23285);
  nand NAND2_4478(II23287,WX6982,II23285);
  nand NAND2_4479(WX7583,II23286,II23287);
  nand NAND2_4480(II23298,WX7062,WX6984);
  nand NAND2_4481(II23299,WX7062,II23298);
  nand NAND2_4482(II23300,WX6984,II23298);
  nand NAND2_4483(WX7590,II23299,II23300);
  nand NAND2_4484(II23311,WX7063,WX6986);
  nand NAND2_4485(II23312,WX7063,II23311);
  nand NAND2_4486(II23313,WX6986,II23311);
  nand NAND2_4487(WX7597,II23312,II23313);
  nand NAND2_4488(II23324,WX7064,WX6988);
  nand NAND2_4489(II23325,WX7064,II23324);
  nand NAND2_4490(II23326,WX6988,II23324);
  nand NAND2_4491(WX7604,II23325,II23326);
  nand NAND2_4492(II23337,WX7065,WX6990);
  nand NAND2_4493(II23338,WX7065,II23337);
  nand NAND2_4494(II23339,WX6990,II23337);
  nand NAND2_4495(WX7611,II23338,II23339);
  nand NAND2_4496(II23350,WX7066,WX6992);
  nand NAND2_4497(II23351,WX7066,II23350);
  nand NAND2_4498(II23352,WX6992,II23350);
  nand NAND2_4499(WX7618,II23351,II23352);
  nand NAND2_4500(II23363,WX7067,WX6994);
  nand NAND2_4501(II23364,WX7067,II23363);
  nand NAND2_4502(II23365,WX6994,II23363);
  nand NAND2_4503(WX7625,II23364,II23365);
  nand NAND2_4504(II23376,WX7068,WX6996);
  nand NAND2_4505(II23377,WX7068,II23376);
  nand NAND2_4506(II23378,WX6996,II23376);
  nand NAND2_4507(WX7632,II23377,II23378);
  nand NAND2_4508(II23389,WX7069,WX6998);
  nand NAND2_4509(II23390,WX7069,II23389);
  nand NAND2_4510(II23391,WX6998,II23389);
  nand NAND2_4511(WX7639,II23390,II23391);
  nand NAND2_4512(II23402,WX7070,WX7000);
  nand NAND2_4513(II23403,WX7070,II23402);
  nand NAND2_4514(II23404,WX7000,II23402);
  nand NAND2_4515(WX7646,II23403,II23404);
  nand NAND2_4516(II23415,WX7071,WX7002);
  nand NAND2_4517(II23416,WX7071,II23415);
  nand NAND2_4518(II23417,WX7002,II23415);
  nand NAND2_4519(WX7653,II23416,II23417);
  nand NAND2_4520(II23428,WX7072,WX7004);
  nand NAND2_4521(II23429,WX7072,II23428);
  nand NAND2_4522(II23430,WX7004,II23428);
  nand NAND2_4523(WX7660,II23429,II23430);
  nand NAND2_4524(II23441,WX7073,WX7006);
  nand NAND2_4525(II23442,WX7073,II23441);
  nand NAND2_4526(II23443,WX7006,II23441);
  nand NAND2_4527(WX7667,II23442,II23443);
  nand NAND2_4528(II23454,WX7074,WX7008);
  nand NAND2_4529(II23455,WX7074,II23454);
  nand NAND2_4530(II23456,WX7008,II23454);
  nand NAND2_4531(WX7674,II23455,II23456);
  nand NAND2_4532(II23467,WX7075,WX7010);
  nand NAND2_4533(II23468,WX7075,II23467);
  nand NAND2_4534(II23469,WX7010,II23467);
  nand NAND2_4535(WX7681,II23468,II23469);
  nand NAND2_4536(II23480,WX7076,WX7012);
  nand NAND2_4537(II23481,WX7076,II23480);
  nand NAND2_4538(II23482,WX7012,II23480);
  nand NAND2_4539(WX7688,II23481,II23482);
  nand NAND2_4540(II23495,WX7092,CRC_OUT_4_31);
  nand NAND2_4541(II23496,WX7092,II23495);
  nand NAND2_4542(II23497,CRC_OUT_4_31,II23495);
  nand NAND2_4543(II23494,II23496,II23497);
  nand NAND2_4544(II23502,CRC_OUT_4_15,II23494);
  nand NAND2_4545(II23503,CRC_OUT_4_15,II23502);
  nand NAND2_4546(II23504,II23494,II23502);
  nand NAND2_4547(WX7696,II23503,II23504);
  nand NAND2_4548(II23510,WX7097,CRC_OUT_4_31);
  nand NAND2_4549(II23511,WX7097,II23510);
  nand NAND2_4550(II23512,CRC_OUT_4_31,II23510);
  nand NAND2_4551(II23509,II23511,II23512);
  nand NAND2_4552(II23517,CRC_OUT_4_10,II23509);
  nand NAND2_4553(II23518,CRC_OUT_4_10,II23517);
  nand NAND2_4554(II23519,II23509,II23517);
  nand NAND2_4555(WX7697,II23518,II23519);
  nand NAND2_4556(II23525,WX7104,CRC_OUT_4_31);
  nand NAND2_4557(II23526,WX7104,II23525);
  nand NAND2_4558(II23527,CRC_OUT_4_31,II23525);
  nand NAND2_4559(II23524,II23526,II23527);
  nand NAND2_4560(II23532,CRC_OUT_4_3,II23524);
  nand NAND2_4561(II23533,CRC_OUT_4_3,II23532);
  nand NAND2_4562(II23534,II23524,II23532);
  nand NAND2_4563(WX7698,II23533,II23534);
  nand NAND2_4564(II23539,WX7108,CRC_OUT_4_31);
  nand NAND2_4565(II23540,WX7108,II23539);
  nand NAND2_4566(II23541,CRC_OUT_4_31,II23539);
  nand NAND2_4567(WX7699,II23540,II23541);
  nand NAND2_4568(II23546,WX7077,CRC_OUT_4_30);
  nand NAND2_4569(II23547,WX7077,II23546);
  nand NAND2_4570(II23548,CRC_OUT_4_30,II23546);
  nand NAND2_4571(WX7700,II23547,II23548);
  nand NAND2_4572(II23553,WX7078,CRC_OUT_4_29);
  nand NAND2_4573(II23554,WX7078,II23553);
  nand NAND2_4574(II23555,CRC_OUT_4_29,II23553);
  nand NAND2_4575(WX7701,II23554,II23555);
  nand NAND2_4576(II23560,WX7079,CRC_OUT_4_28);
  nand NAND2_4577(II23561,WX7079,II23560);
  nand NAND2_4578(II23562,CRC_OUT_4_28,II23560);
  nand NAND2_4579(WX7702,II23561,II23562);
  nand NAND2_4580(II23567,WX7080,CRC_OUT_4_27);
  nand NAND2_4581(II23568,WX7080,II23567);
  nand NAND2_4582(II23569,CRC_OUT_4_27,II23567);
  nand NAND2_4583(WX7703,II23568,II23569);
  nand NAND2_4584(II23574,WX7081,CRC_OUT_4_26);
  nand NAND2_4585(II23575,WX7081,II23574);
  nand NAND2_4586(II23576,CRC_OUT_4_26,II23574);
  nand NAND2_4587(WX7704,II23575,II23576);
  nand NAND2_4588(II23581,WX7082,CRC_OUT_4_25);
  nand NAND2_4589(II23582,WX7082,II23581);
  nand NAND2_4590(II23583,CRC_OUT_4_25,II23581);
  nand NAND2_4591(WX7705,II23582,II23583);
  nand NAND2_4592(II23588,WX7083,CRC_OUT_4_24);
  nand NAND2_4593(II23589,WX7083,II23588);
  nand NAND2_4594(II23590,CRC_OUT_4_24,II23588);
  nand NAND2_4595(WX7706,II23589,II23590);
  nand NAND2_4596(II23595,WX7084,CRC_OUT_4_23);
  nand NAND2_4597(II23596,WX7084,II23595);
  nand NAND2_4598(II23597,CRC_OUT_4_23,II23595);
  nand NAND2_4599(WX7707,II23596,II23597);
  nand NAND2_4600(II23602,WX7085,CRC_OUT_4_22);
  nand NAND2_4601(II23603,WX7085,II23602);
  nand NAND2_4602(II23604,CRC_OUT_4_22,II23602);
  nand NAND2_4603(WX7708,II23603,II23604);
  nand NAND2_4604(II23609,WX7086,CRC_OUT_4_21);
  nand NAND2_4605(II23610,WX7086,II23609);
  nand NAND2_4606(II23611,CRC_OUT_4_21,II23609);
  nand NAND2_4607(WX7709,II23610,II23611);
  nand NAND2_4608(II23616,WX7087,CRC_OUT_4_20);
  nand NAND2_4609(II23617,WX7087,II23616);
  nand NAND2_4610(II23618,CRC_OUT_4_20,II23616);
  nand NAND2_4611(WX7710,II23617,II23618);
  nand NAND2_4612(II23623,WX7088,CRC_OUT_4_19);
  nand NAND2_4613(II23624,WX7088,II23623);
  nand NAND2_4614(II23625,CRC_OUT_4_19,II23623);
  nand NAND2_4615(WX7711,II23624,II23625);
  nand NAND2_4616(II23630,WX7089,CRC_OUT_4_18);
  nand NAND2_4617(II23631,WX7089,II23630);
  nand NAND2_4618(II23632,CRC_OUT_4_18,II23630);
  nand NAND2_4619(WX7712,II23631,II23632);
  nand NAND2_4620(II23637,WX7090,CRC_OUT_4_17);
  nand NAND2_4621(II23638,WX7090,II23637);
  nand NAND2_4622(II23639,CRC_OUT_4_17,II23637);
  nand NAND2_4623(WX7713,II23638,II23639);
  nand NAND2_4624(II23644,WX7091,CRC_OUT_4_16);
  nand NAND2_4625(II23645,WX7091,II23644);
  nand NAND2_4626(II23646,CRC_OUT_4_16,II23644);
  nand NAND2_4627(WX7714,II23645,II23646);
  nand NAND2_4628(II23651,WX7093,CRC_OUT_4_14);
  nand NAND2_4629(II23652,WX7093,II23651);
  nand NAND2_4630(II23653,CRC_OUT_4_14,II23651);
  nand NAND2_4631(WX7715,II23652,II23653);
  nand NAND2_4632(II23658,WX7094,CRC_OUT_4_13);
  nand NAND2_4633(II23659,WX7094,II23658);
  nand NAND2_4634(II23660,CRC_OUT_4_13,II23658);
  nand NAND2_4635(WX7716,II23659,II23660);
  nand NAND2_4636(II23665,WX7095,CRC_OUT_4_12);
  nand NAND2_4637(II23666,WX7095,II23665);
  nand NAND2_4638(II23667,CRC_OUT_4_12,II23665);
  nand NAND2_4639(WX7717,II23666,II23667);
  nand NAND2_4640(II23672,WX7096,CRC_OUT_4_11);
  nand NAND2_4641(II23673,WX7096,II23672);
  nand NAND2_4642(II23674,CRC_OUT_4_11,II23672);
  nand NAND2_4643(WX7718,II23673,II23674);
  nand NAND2_4644(II23679,WX7098,CRC_OUT_4_9);
  nand NAND2_4645(II23680,WX7098,II23679);
  nand NAND2_4646(II23681,CRC_OUT_4_9,II23679);
  nand NAND2_4647(WX7719,II23680,II23681);
  nand NAND2_4648(II23686,WX7099,CRC_OUT_4_8);
  nand NAND2_4649(II23687,WX7099,II23686);
  nand NAND2_4650(II23688,CRC_OUT_4_8,II23686);
  nand NAND2_4651(WX7720,II23687,II23688);
  nand NAND2_4652(II23693,WX7100,CRC_OUT_4_7);
  nand NAND2_4653(II23694,WX7100,II23693);
  nand NAND2_4654(II23695,CRC_OUT_4_7,II23693);
  nand NAND2_4655(WX7721,II23694,II23695);
  nand NAND2_4656(II23700,WX7101,CRC_OUT_4_6);
  nand NAND2_4657(II23701,WX7101,II23700);
  nand NAND2_4658(II23702,CRC_OUT_4_6,II23700);
  nand NAND2_4659(WX7722,II23701,II23702);
  nand NAND2_4660(II23707,WX7102,CRC_OUT_4_5);
  nand NAND2_4661(II23708,WX7102,II23707);
  nand NAND2_4662(II23709,CRC_OUT_4_5,II23707);
  nand NAND2_4663(WX7723,II23708,II23709);
  nand NAND2_4664(II23714,WX7103,CRC_OUT_4_4);
  nand NAND2_4665(II23715,WX7103,II23714);
  nand NAND2_4666(II23716,CRC_OUT_4_4,II23714);
  nand NAND2_4667(WX7724,II23715,II23716);
  nand NAND2_4668(II23721,WX7105,CRC_OUT_4_2);
  nand NAND2_4669(II23722,WX7105,II23721);
  nand NAND2_4670(II23723,CRC_OUT_4_2,II23721);
  nand NAND2_4671(WX7725,II23722,II23723);
  nand NAND2_4672(II23728,WX7106,CRC_OUT_4_1);
  nand NAND2_4673(II23729,WX7106,II23728);
  nand NAND2_4674(II23730,CRC_OUT_4_1,II23728);
  nand NAND2_4675(WX7726,II23729,II23730);
  nand NAND2_4676(II23735,WX7107,CRC_OUT_4_0);
  nand NAND2_4677(II23736,WX7107,II23735);
  nand NAND2_4678(II23737,CRC_OUT_4_0,II23735);
  nand NAND2_4679(WX7727,II23736,II23737);
  nand NAND2_4680(II26018,WX8759,WX8403);
  nand NAND2_4681(II26019,WX8759,II26018);
  nand NAND2_4682(II26020,WX8403,II26018);
  nand NAND2_4683(II26017,II26019,II26020);
  nand NAND2_4684(II26025,WX8467,II26017);
  nand NAND2_4685(II26026,WX8467,II26025);
  nand NAND2_4686(II26027,II26017,II26025);
  nand NAND2_4687(II26016,II26026,II26027);
  nand NAND2_4688(II26033,WX8531,WX8595);
  nand NAND2_4689(II26034,WX8531,II26033);
  nand NAND2_4690(II26035,WX8595,II26033);
  nand NAND2_4691(II26032,II26034,II26035);
  nand NAND2_4692(II26040,II26016,II26032);
  nand NAND2_4693(II26041,II26016,II26040);
  nand NAND2_4694(II26042,II26032,II26040);
  nand NAND2_4695(WX8658,II26041,II26042);
  nand NAND2_4696(II26049,WX8759,WX8405);
  nand NAND2_4697(II26050,WX8759,II26049);
  nand NAND2_4698(II26051,WX8405,II26049);
  nand NAND2_4699(II26048,II26050,II26051);
  nand NAND2_4700(II26056,WX8469,II26048);
  nand NAND2_4701(II26057,WX8469,II26056);
  nand NAND2_4702(II26058,II26048,II26056);
  nand NAND2_4703(II26047,II26057,II26058);
  nand NAND2_4704(II26064,WX8533,WX8597);
  nand NAND2_4705(II26065,WX8533,II26064);
  nand NAND2_4706(II26066,WX8597,II26064);
  nand NAND2_4707(II26063,II26065,II26066);
  nand NAND2_4708(II26071,II26047,II26063);
  nand NAND2_4709(II26072,II26047,II26071);
  nand NAND2_4710(II26073,II26063,II26071);
  nand NAND2_4711(WX8659,II26072,II26073);
  nand NAND2_4712(II26080,WX8759,WX8407);
  nand NAND2_4713(II26081,WX8759,II26080);
  nand NAND2_4714(II26082,WX8407,II26080);
  nand NAND2_4715(II26079,II26081,II26082);
  nand NAND2_4716(II26087,WX8471,II26079);
  nand NAND2_4717(II26088,WX8471,II26087);
  nand NAND2_4718(II26089,II26079,II26087);
  nand NAND2_4719(II26078,II26088,II26089);
  nand NAND2_4720(II26095,WX8535,WX8599);
  nand NAND2_4721(II26096,WX8535,II26095);
  nand NAND2_4722(II26097,WX8599,II26095);
  nand NAND2_4723(II26094,II26096,II26097);
  nand NAND2_4724(II26102,II26078,II26094);
  nand NAND2_4725(II26103,II26078,II26102);
  nand NAND2_4726(II26104,II26094,II26102);
  nand NAND2_4727(WX8660,II26103,II26104);
  nand NAND2_4728(II26111,WX8759,WX8409);
  nand NAND2_4729(II26112,WX8759,II26111);
  nand NAND2_4730(II26113,WX8409,II26111);
  nand NAND2_4731(II26110,II26112,II26113);
  nand NAND2_4732(II26118,WX8473,II26110);
  nand NAND2_4733(II26119,WX8473,II26118);
  nand NAND2_4734(II26120,II26110,II26118);
  nand NAND2_4735(II26109,II26119,II26120);
  nand NAND2_4736(II26126,WX8537,WX8601);
  nand NAND2_4737(II26127,WX8537,II26126);
  nand NAND2_4738(II26128,WX8601,II26126);
  nand NAND2_4739(II26125,II26127,II26128);
  nand NAND2_4740(II26133,II26109,II26125);
  nand NAND2_4741(II26134,II26109,II26133);
  nand NAND2_4742(II26135,II26125,II26133);
  nand NAND2_4743(WX8661,II26134,II26135);
  nand NAND2_4744(II26142,WX8759,WX8411);
  nand NAND2_4745(II26143,WX8759,II26142);
  nand NAND2_4746(II26144,WX8411,II26142);
  nand NAND2_4747(II26141,II26143,II26144);
  nand NAND2_4748(II26149,WX8475,II26141);
  nand NAND2_4749(II26150,WX8475,II26149);
  nand NAND2_4750(II26151,II26141,II26149);
  nand NAND2_4751(II26140,II26150,II26151);
  nand NAND2_4752(II26157,WX8539,WX8603);
  nand NAND2_4753(II26158,WX8539,II26157);
  nand NAND2_4754(II26159,WX8603,II26157);
  nand NAND2_4755(II26156,II26158,II26159);
  nand NAND2_4756(II26164,II26140,II26156);
  nand NAND2_4757(II26165,II26140,II26164);
  nand NAND2_4758(II26166,II26156,II26164);
  nand NAND2_4759(WX8662,II26165,II26166);
  nand NAND2_4760(II26173,WX8759,WX8413);
  nand NAND2_4761(II26174,WX8759,II26173);
  nand NAND2_4762(II26175,WX8413,II26173);
  nand NAND2_4763(II26172,II26174,II26175);
  nand NAND2_4764(II26180,WX8477,II26172);
  nand NAND2_4765(II26181,WX8477,II26180);
  nand NAND2_4766(II26182,II26172,II26180);
  nand NAND2_4767(II26171,II26181,II26182);
  nand NAND2_4768(II26188,WX8541,WX8605);
  nand NAND2_4769(II26189,WX8541,II26188);
  nand NAND2_4770(II26190,WX8605,II26188);
  nand NAND2_4771(II26187,II26189,II26190);
  nand NAND2_4772(II26195,II26171,II26187);
  nand NAND2_4773(II26196,II26171,II26195);
  nand NAND2_4774(II26197,II26187,II26195);
  nand NAND2_4775(WX8663,II26196,II26197);
  nand NAND2_4776(II26204,WX8759,WX8415);
  nand NAND2_4777(II26205,WX8759,II26204);
  nand NAND2_4778(II26206,WX8415,II26204);
  nand NAND2_4779(II26203,II26205,II26206);
  nand NAND2_4780(II26211,WX8479,II26203);
  nand NAND2_4781(II26212,WX8479,II26211);
  nand NAND2_4782(II26213,II26203,II26211);
  nand NAND2_4783(II26202,II26212,II26213);
  nand NAND2_4784(II26219,WX8543,WX8607);
  nand NAND2_4785(II26220,WX8543,II26219);
  nand NAND2_4786(II26221,WX8607,II26219);
  nand NAND2_4787(II26218,II26220,II26221);
  nand NAND2_4788(II26226,II26202,II26218);
  nand NAND2_4789(II26227,II26202,II26226);
  nand NAND2_4790(II26228,II26218,II26226);
  nand NAND2_4791(WX8664,II26227,II26228);
  nand NAND2_4792(II26235,WX8759,WX8417);
  nand NAND2_4793(II26236,WX8759,II26235);
  nand NAND2_4794(II26237,WX8417,II26235);
  nand NAND2_4795(II26234,II26236,II26237);
  nand NAND2_4796(II26242,WX8481,II26234);
  nand NAND2_4797(II26243,WX8481,II26242);
  nand NAND2_4798(II26244,II26234,II26242);
  nand NAND2_4799(II26233,II26243,II26244);
  nand NAND2_4800(II26250,WX8545,WX8609);
  nand NAND2_4801(II26251,WX8545,II26250);
  nand NAND2_4802(II26252,WX8609,II26250);
  nand NAND2_4803(II26249,II26251,II26252);
  nand NAND2_4804(II26257,II26233,II26249);
  nand NAND2_4805(II26258,II26233,II26257);
  nand NAND2_4806(II26259,II26249,II26257);
  nand NAND2_4807(WX8665,II26258,II26259);
  nand NAND2_4808(II26266,WX8759,WX8419);
  nand NAND2_4809(II26267,WX8759,II26266);
  nand NAND2_4810(II26268,WX8419,II26266);
  nand NAND2_4811(II26265,II26267,II26268);
  nand NAND2_4812(II26273,WX8483,II26265);
  nand NAND2_4813(II26274,WX8483,II26273);
  nand NAND2_4814(II26275,II26265,II26273);
  nand NAND2_4815(II26264,II26274,II26275);
  nand NAND2_4816(II26281,WX8547,WX8611);
  nand NAND2_4817(II26282,WX8547,II26281);
  nand NAND2_4818(II26283,WX8611,II26281);
  nand NAND2_4819(II26280,II26282,II26283);
  nand NAND2_4820(II26288,II26264,II26280);
  nand NAND2_4821(II26289,II26264,II26288);
  nand NAND2_4822(II26290,II26280,II26288);
  nand NAND2_4823(WX8666,II26289,II26290);
  nand NAND2_4824(II26297,WX8759,WX8421);
  nand NAND2_4825(II26298,WX8759,II26297);
  nand NAND2_4826(II26299,WX8421,II26297);
  nand NAND2_4827(II26296,II26298,II26299);
  nand NAND2_4828(II26304,WX8485,II26296);
  nand NAND2_4829(II26305,WX8485,II26304);
  nand NAND2_4830(II26306,II26296,II26304);
  nand NAND2_4831(II26295,II26305,II26306);
  nand NAND2_4832(II26312,WX8549,WX8613);
  nand NAND2_4833(II26313,WX8549,II26312);
  nand NAND2_4834(II26314,WX8613,II26312);
  nand NAND2_4835(II26311,II26313,II26314);
  nand NAND2_4836(II26319,II26295,II26311);
  nand NAND2_4837(II26320,II26295,II26319);
  nand NAND2_4838(II26321,II26311,II26319);
  nand NAND2_4839(WX8667,II26320,II26321);
  nand NAND2_4840(II26328,WX8759,WX8423);
  nand NAND2_4841(II26329,WX8759,II26328);
  nand NAND2_4842(II26330,WX8423,II26328);
  nand NAND2_4843(II26327,II26329,II26330);
  nand NAND2_4844(II26335,WX8487,II26327);
  nand NAND2_4845(II26336,WX8487,II26335);
  nand NAND2_4846(II26337,II26327,II26335);
  nand NAND2_4847(II26326,II26336,II26337);
  nand NAND2_4848(II26343,WX8551,WX8615);
  nand NAND2_4849(II26344,WX8551,II26343);
  nand NAND2_4850(II26345,WX8615,II26343);
  nand NAND2_4851(II26342,II26344,II26345);
  nand NAND2_4852(II26350,II26326,II26342);
  nand NAND2_4853(II26351,II26326,II26350);
  nand NAND2_4854(II26352,II26342,II26350);
  nand NAND2_4855(WX8668,II26351,II26352);
  nand NAND2_4856(II26359,WX8759,WX8425);
  nand NAND2_4857(II26360,WX8759,II26359);
  nand NAND2_4858(II26361,WX8425,II26359);
  nand NAND2_4859(II26358,II26360,II26361);
  nand NAND2_4860(II26366,WX8489,II26358);
  nand NAND2_4861(II26367,WX8489,II26366);
  nand NAND2_4862(II26368,II26358,II26366);
  nand NAND2_4863(II26357,II26367,II26368);
  nand NAND2_4864(II26374,WX8553,WX8617);
  nand NAND2_4865(II26375,WX8553,II26374);
  nand NAND2_4866(II26376,WX8617,II26374);
  nand NAND2_4867(II26373,II26375,II26376);
  nand NAND2_4868(II26381,II26357,II26373);
  nand NAND2_4869(II26382,II26357,II26381);
  nand NAND2_4870(II26383,II26373,II26381);
  nand NAND2_4871(WX8669,II26382,II26383);
  nand NAND2_4872(II26390,WX8759,WX8427);
  nand NAND2_4873(II26391,WX8759,II26390);
  nand NAND2_4874(II26392,WX8427,II26390);
  nand NAND2_4875(II26389,II26391,II26392);
  nand NAND2_4876(II26397,WX8491,II26389);
  nand NAND2_4877(II26398,WX8491,II26397);
  nand NAND2_4878(II26399,II26389,II26397);
  nand NAND2_4879(II26388,II26398,II26399);
  nand NAND2_4880(II26405,WX8555,WX8619);
  nand NAND2_4881(II26406,WX8555,II26405);
  nand NAND2_4882(II26407,WX8619,II26405);
  nand NAND2_4883(II26404,II26406,II26407);
  nand NAND2_4884(II26412,II26388,II26404);
  nand NAND2_4885(II26413,II26388,II26412);
  nand NAND2_4886(II26414,II26404,II26412);
  nand NAND2_4887(WX8670,II26413,II26414);
  nand NAND2_4888(II26421,WX8759,WX8429);
  nand NAND2_4889(II26422,WX8759,II26421);
  nand NAND2_4890(II26423,WX8429,II26421);
  nand NAND2_4891(II26420,II26422,II26423);
  nand NAND2_4892(II26428,WX8493,II26420);
  nand NAND2_4893(II26429,WX8493,II26428);
  nand NAND2_4894(II26430,II26420,II26428);
  nand NAND2_4895(II26419,II26429,II26430);
  nand NAND2_4896(II26436,WX8557,WX8621);
  nand NAND2_4897(II26437,WX8557,II26436);
  nand NAND2_4898(II26438,WX8621,II26436);
  nand NAND2_4899(II26435,II26437,II26438);
  nand NAND2_4900(II26443,II26419,II26435);
  nand NAND2_4901(II26444,II26419,II26443);
  nand NAND2_4902(II26445,II26435,II26443);
  nand NAND2_4903(WX8671,II26444,II26445);
  nand NAND2_4904(II26452,WX8759,WX8431);
  nand NAND2_4905(II26453,WX8759,II26452);
  nand NAND2_4906(II26454,WX8431,II26452);
  nand NAND2_4907(II26451,II26453,II26454);
  nand NAND2_4908(II26459,WX8495,II26451);
  nand NAND2_4909(II26460,WX8495,II26459);
  nand NAND2_4910(II26461,II26451,II26459);
  nand NAND2_4911(II26450,II26460,II26461);
  nand NAND2_4912(II26467,WX8559,WX8623);
  nand NAND2_4913(II26468,WX8559,II26467);
  nand NAND2_4914(II26469,WX8623,II26467);
  nand NAND2_4915(II26466,II26468,II26469);
  nand NAND2_4916(II26474,II26450,II26466);
  nand NAND2_4917(II26475,II26450,II26474);
  nand NAND2_4918(II26476,II26466,II26474);
  nand NAND2_4919(WX8672,II26475,II26476);
  nand NAND2_4920(II26483,WX8759,WX8433);
  nand NAND2_4921(II26484,WX8759,II26483);
  nand NAND2_4922(II26485,WX8433,II26483);
  nand NAND2_4923(II26482,II26484,II26485);
  nand NAND2_4924(II26490,WX8497,II26482);
  nand NAND2_4925(II26491,WX8497,II26490);
  nand NAND2_4926(II26492,II26482,II26490);
  nand NAND2_4927(II26481,II26491,II26492);
  nand NAND2_4928(II26498,WX8561,WX8625);
  nand NAND2_4929(II26499,WX8561,II26498);
  nand NAND2_4930(II26500,WX8625,II26498);
  nand NAND2_4931(II26497,II26499,II26500);
  nand NAND2_4932(II26505,II26481,II26497);
  nand NAND2_4933(II26506,II26481,II26505);
  nand NAND2_4934(II26507,II26497,II26505);
  nand NAND2_4935(WX8673,II26506,II26507);
  nand NAND2_4936(II26514,WX8760,WX8435);
  nand NAND2_4937(II26515,WX8760,II26514);
  nand NAND2_4938(II26516,WX8435,II26514);
  nand NAND2_4939(II26513,II26515,II26516);
  nand NAND2_4940(II26521,WX8499,II26513);
  nand NAND2_4941(II26522,WX8499,II26521);
  nand NAND2_4942(II26523,II26513,II26521);
  nand NAND2_4943(II26512,II26522,II26523);
  nand NAND2_4944(II26529,WX8563,WX8627);
  nand NAND2_4945(II26530,WX8563,II26529);
  nand NAND2_4946(II26531,WX8627,II26529);
  nand NAND2_4947(II26528,II26530,II26531);
  nand NAND2_4948(II26536,II26512,II26528);
  nand NAND2_4949(II26537,II26512,II26536);
  nand NAND2_4950(II26538,II26528,II26536);
  nand NAND2_4951(WX8674,II26537,II26538);
  nand NAND2_4952(II26545,WX8760,WX8437);
  nand NAND2_4953(II26546,WX8760,II26545);
  nand NAND2_4954(II26547,WX8437,II26545);
  nand NAND2_4955(II26544,II26546,II26547);
  nand NAND2_4956(II26552,WX8501,II26544);
  nand NAND2_4957(II26553,WX8501,II26552);
  nand NAND2_4958(II26554,II26544,II26552);
  nand NAND2_4959(II26543,II26553,II26554);
  nand NAND2_4960(II26560,WX8565,WX8629);
  nand NAND2_4961(II26561,WX8565,II26560);
  nand NAND2_4962(II26562,WX8629,II26560);
  nand NAND2_4963(II26559,II26561,II26562);
  nand NAND2_4964(II26567,II26543,II26559);
  nand NAND2_4965(II26568,II26543,II26567);
  nand NAND2_4966(II26569,II26559,II26567);
  nand NAND2_4967(WX8675,II26568,II26569);
  nand NAND2_4968(II26576,WX8760,WX8439);
  nand NAND2_4969(II26577,WX8760,II26576);
  nand NAND2_4970(II26578,WX8439,II26576);
  nand NAND2_4971(II26575,II26577,II26578);
  nand NAND2_4972(II26583,WX8503,II26575);
  nand NAND2_4973(II26584,WX8503,II26583);
  nand NAND2_4974(II26585,II26575,II26583);
  nand NAND2_4975(II26574,II26584,II26585);
  nand NAND2_4976(II26591,WX8567,WX8631);
  nand NAND2_4977(II26592,WX8567,II26591);
  nand NAND2_4978(II26593,WX8631,II26591);
  nand NAND2_4979(II26590,II26592,II26593);
  nand NAND2_4980(II26598,II26574,II26590);
  nand NAND2_4981(II26599,II26574,II26598);
  nand NAND2_4982(II26600,II26590,II26598);
  nand NAND2_4983(WX8676,II26599,II26600);
  nand NAND2_4984(II26607,WX8760,WX8441);
  nand NAND2_4985(II26608,WX8760,II26607);
  nand NAND2_4986(II26609,WX8441,II26607);
  nand NAND2_4987(II26606,II26608,II26609);
  nand NAND2_4988(II26614,WX8505,II26606);
  nand NAND2_4989(II26615,WX8505,II26614);
  nand NAND2_4990(II26616,II26606,II26614);
  nand NAND2_4991(II26605,II26615,II26616);
  nand NAND2_4992(II26622,WX8569,WX8633);
  nand NAND2_4993(II26623,WX8569,II26622);
  nand NAND2_4994(II26624,WX8633,II26622);
  nand NAND2_4995(II26621,II26623,II26624);
  nand NAND2_4996(II26629,II26605,II26621);
  nand NAND2_4997(II26630,II26605,II26629);
  nand NAND2_4998(II26631,II26621,II26629);
  nand NAND2_4999(WX8677,II26630,II26631);
  nand NAND2_5000(II26638,WX8760,WX8443);
  nand NAND2_5001(II26639,WX8760,II26638);
  nand NAND2_5002(II26640,WX8443,II26638);
  nand NAND2_5003(II26637,II26639,II26640);
  nand NAND2_5004(II26645,WX8507,II26637);
  nand NAND2_5005(II26646,WX8507,II26645);
  nand NAND2_5006(II26647,II26637,II26645);
  nand NAND2_5007(II26636,II26646,II26647);
  nand NAND2_5008(II26653,WX8571,WX8635);
  nand NAND2_5009(II26654,WX8571,II26653);
  nand NAND2_5010(II26655,WX8635,II26653);
  nand NAND2_5011(II26652,II26654,II26655);
  nand NAND2_5012(II26660,II26636,II26652);
  nand NAND2_5013(II26661,II26636,II26660);
  nand NAND2_5014(II26662,II26652,II26660);
  nand NAND2_5015(WX8678,II26661,II26662);
  nand NAND2_5016(II26669,WX8760,WX8445);
  nand NAND2_5017(II26670,WX8760,II26669);
  nand NAND2_5018(II26671,WX8445,II26669);
  nand NAND2_5019(II26668,II26670,II26671);
  nand NAND2_5020(II26676,WX8509,II26668);
  nand NAND2_5021(II26677,WX8509,II26676);
  nand NAND2_5022(II26678,II26668,II26676);
  nand NAND2_5023(II26667,II26677,II26678);
  nand NAND2_5024(II26684,WX8573,WX8637);
  nand NAND2_5025(II26685,WX8573,II26684);
  nand NAND2_5026(II26686,WX8637,II26684);
  nand NAND2_5027(II26683,II26685,II26686);
  nand NAND2_5028(II26691,II26667,II26683);
  nand NAND2_5029(II26692,II26667,II26691);
  nand NAND2_5030(II26693,II26683,II26691);
  nand NAND2_5031(WX8679,II26692,II26693);
  nand NAND2_5032(II26700,WX8760,WX8447);
  nand NAND2_5033(II26701,WX8760,II26700);
  nand NAND2_5034(II26702,WX8447,II26700);
  nand NAND2_5035(II26699,II26701,II26702);
  nand NAND2_5036(II26707,WX8511,II26699);
  nand NAND2_5037(II26708,WX8511,II26707);
  nand NAND2_5038(II26709,II26699,II26707);
  nand NAND2_5039(II26698,II26708,II26709);
  nand NAND2_5040(II26715,WX8575,WX8639);
  nand NAND2_5041(II26716,WX8575,II26715);
  nand NAND2_5042(II26717,WX8639,II26715);
  nand NAND2_5043(II26714,II26716,II26717);
  nand NAND2_5044(II26722,II26698,II26714);
  nand NAND2_5045(II26723,II26698,II26722);
  nand NAND2_5046(II26724,II26714,II26722);
  nand NAND2_5047(WX8680,II26723,II26724);
  nand NAND2_5048(II26731,WX8760,WX8449);
  nand NAND2_5049(II26732,WX8760,II26731);
  nand NAND2_5050(II26733,WX8449,II26731);
  nand NAND2_5051(II26730,II26732,II26733);
  nand NAND2_5052(II26738,WX8513,II26730);
  nand NAND2_5053(II26739,WX8513,II26738);
  nand NAND2_5054(II26740,II26730,II26738);
  nand NAND2_5055(II26729,II26739,II26740);
  nand NAND2_5056(II26746,WX8577,WX8641);
  nand NAND2_5057(II26747,WX8577,II26746);
  nand NAND2_5058(II26748,WX8641,II26746);
  nand NAND2_5059(II26745,II26747,II26748);
  nand NAND2_5060(II26753,II26729,II26745);
  nand NAND2_5061(II26754,II26729,II26753);
  nand NAND2_5062(II26755,II26745,II26753);
  nand NAND2_5063(WX8681,II26754,II26755);
  nand NAND2_5064(II26762,WX8760,WX8451);
  nand NAND2_5065(II26763,WX8760,II26762);
  nand NAND2_5066(II26764,WX8451,II26762);
  nand NAND2_5067(II26761,II26763,II26764);
  nand NAND2_5068(II26769,WX8515,II26761);
  nand NAND2_5069(II26770,WX8515,II26769);
  nand NAND2_5070(II26771,II26761,II26769);
  nand NAND2_5071(II26760,II26770,II26771);
  nand NAND2_5072(II26777,WX8579,WX8643);
  nand NAND2_5073(II26778,WX8579,II26777);
  nand NAND2_5074(II26779,WX8643,II26777);
  nand NAND2_5075(II26776,II26778,II26779);
  nand NAND2_5076(II26784,II26760,II26776);
  nand NAND2_5077(II26785,II26760,II26784);
  nand NAND2_5078(II26786,II26776,II26784);
  nand NAND2_5079(WX8682,II26785,II26786);
  nand NAND2_5080(II26793,WX8760,WX8453);
  nand NAND2_5081(II26794,WX8760,II26793);
  nand NAND2_5082(II26795,WX8453,II26793);
  nand NAND2_5083(II26792,II26794,II26795);
  nand NAND2_5084(II26800,WX8517,II26792);
  nand NAND2_5085(II26801,WX8517,II26800);
  nand NAND2_5086(II26802,II26792,II26800);
  nand NAND2_5087(II26791,II26801,II26802);
  nand NAND2_5088(II26808,WX8581,WX8645);
  nand NAND2_5089(II26809,WX8581,II26808);
  nand NAND2_5090(II26810,WX8645,II26808);
  nand NAND2_5091(II26807,II26809,II26810);
  nand NAND2_5092(II26815,II26791,II26807);
  nand NAND2_5093(II26816,II26791,II26815);
  nand NAND2_5094(II26817,II26807,II26815);
  nand NAND2_5095(WX8683,II26816,II26817);
  nand NAND2_5096(II26824,WX8760,WX8455);
  nand NAND2_5097(II26825,WX8760,II26824);
  nand NAND2_5098(II26826,WX8455,II26824);
  nand NAND2_5099(II26823,II26825,II26826);
  nand NAND2_5100(II26831,WX8519,II26823);
  nand NAND2_5101(II26832,WX8519,II26831);
  nand NAND2_5102(II26833,II26823,II26831);
  nand NAND2_5103(II26822,II26832,II26833);
  nand NAND2_5104(II26839,WX8583,WX8647);
  nand NAND2_5105(II26840,WX8583,II26839);
  nand NAND2_5106(II26841,WX8647,II26839);
  nand NAND2_5107(II26838,II26840,II26841);
  nand NAND2_5108(II26846,II26822,II26838);
  nand NAND2_5109(II26847,II26822,II26846);
  nand NAND2_5110(II26848,II26838,II26846);
  nand NAND2_5111(WX8684,II26847,II26848);
  nand NAND2_5112(II26855,WX8760,WX8457);
  nand NAND2_5113(II26856,WX8760,II26855);
  nand NAND2_5114(II26857,WX8457,II26855);
  nand NAND2_5115(II26854,II26856,II26857);
  nand NAND2_5116(II26862,WX8521,II26854);
  nand NAND2_5117(II26863,WX8521,II26862);
  nand NAND2_5118(II26864,II26854,II26862);
  nand NAND2_5119(II26853,II26863,II26864);
  nand NAND2_5120(II26870,WX8585,WX8649);
  nand NAND2_5121(II26871,WX8585,II26870);
  nand NAND2_5122(II26872,WX8649,II26870);
  nand NAND2_5123(II26869,II26871,II26872);
  nand NAND2_5124(II26877,II26853,II26869);
  nand NAND2_5125(II26878,II26853,II26877);
  nand NAND2_5126(II26879,II26869,II26877);
  nand NAND2_5127(WX8685,II26878,II26879);
  nand NAND2_5128(II26886,WX8760,WX8459);
  nand NAND2_5129(II26887,WX8760,II26886);
  nand NAND2_5130(II26888,WX8459,II26886);
  nand NAND2_5131(II26885,II26887,II26888);
  nand NAND2_5132(II26893,WX8523,II26885);
  nand NAND2_5133(II26894,WX8523,II26893);
  nand NAND2_5134(II26895,II26885,II26893);
  nand NAND2_5135(II26884,II26894,II26895);
  nand NAND2_5136(II26901,WX8587,WX8651);
  nand NAND2_5137(II26902,WX8587,II26901);
  nand NAND2_5138(II26903,WX8651,II26901);
  nand NAND2_5139(II26900,II26902,II26903);
  nand NAND2_5140(II26908,II26884,II26900);
  nand NAND2_5141(II26909,II26884,II26908);
  nand NAND2_5142(II26910,II26900,II26908);
  nand NAND2_5143(WX8686,II26909,II26910);
  nand NAND2_5144(II26917,WX8760,WX8461);
  nand NAND2_5145(II26918,WX8760,II26917);
  nand NAND2_5146(II26919,WX8461,II26917);
  nand NAND2_5147(II26916,II26918,II26919);
  nand NAND2_5148(II26924,WX8525,II26916);
  nand NAND2_5149(II26925,WX8525,II26924);
  nand NAND2_5150(II26926,II26916,II26924);
  nand NAND2_5151(II26915,II26925,II26926);
  nand NAND2_5152(II26932,WX8589,WX8653);
  nand NAND2_5153(II26933,WX8589,II26932);
  nand NAND2_5154(II26934,WX8653,II26932);
  nand NAND2_5155(II26931,II26933,II26934);
  nand NAND2_5156(II26939,II26915,II26931);
  nand NAND2_5157(II26940,II26915,II26939);
  nand NAND2_5158(II26941,II26931,II26939);
  nand NAND2_5159(WX8687,II26940,II26941);
  nand NAND2_5160(II26948,WX8760,WX8463);
  nand NAND2_5161(II26949,WX8760,II26948);
  nand NAND2_5162(II26950,WX8463,II26948);
  nand NAND2_5163(II26947,II26949,II26950);
  nand NAND2_5164(II26955,WX8527,II26947);
  nand NAND2_5165(II26956,WX8527,II26955);
  nand NAND2_5166(II26957,II26947,II26955);
  nand NAND2_5167(II26946,II26956,II26957);
  nand NAND2_5168(II26963,WX8591,WX8655);
  nand NAND2_5169(II26964,WX8591,II26963);
  nand NAND2_5170(II26965,WX8655,II26963);
  nand NAND2_5171(II26962,II26964,II26965);
  nand NAND2_5172(II26970,II26946,II26962);
  nand NAND2_5173(II26971,II26946,II26970);
  nand NAND2_5174(II26972,II26962,II26970);
  nand NAND2_5175(WX8688,II26971,II26972);
  nand NAND2_5176(II26979,WX8760,WX8465);
  nand NAND2_5177(II26980,WX8760,II26979);
  nand NAND2_5178(II26981,WX8465,II26979);
  nand NAND2_5179(II26978,II26980,II26981);
  nand NAND2_5180(II26986,WX8529,II26978);
  nand NAND2_5181(II26987,WX8529,II26986);
  nand NAND2_5182(II26988,II26978,II26986);
  nand NAND2_5183(II26977,II26987,II26988);
  nand NAND2_5184(II26994,WX8593,WX8657);
  nand NAND2_5185(II26995,WX8593,II26994);
  nand NAND2_5186(II26996,WX8657,II26994);
  nand NAND2_5187(II26993,II26995,II26996);
  nand NAND2_5188(II27001,II26977,II26993);
  nand NAND2_5189(II27002,II26977,II27001);
  nand NAND2_5190(II27003,II26993,II27001);
  nand NAND2_5191(WX8689,II27002,II27003);
  nand NAND2_5192(II27082,WX8338,WX8243);
  nand NAND2_5193(II27083,WX8338,II27082);
  nand NAND2_5194(II27084,WX8243,II27082);
  nand NAND2_5195(WX8764,II27083,II27084);
  nand NAND2_5196(II27095,WX8339,WX8245);
  nand NAND2_5197(II27096,WX8339,II27095);
  nand NAND2_5198(II27097,WX8245,II27095);
  nand NAND2_5199(WX8771,II27096,II27097);
  nand NAND2_5200(II27108,WX8340,WX8247);
  nand NAND2_5201(II27109,WX8340,II27108);
  nand NAND2_5202(II27110,WX8247,II27108);
  nand NAND2_5203(WX8778,II27109,II27110);
  nand NAND2_5204(II27121,WX8341,WX8249);
  nand NAND2_5205(II27122,WX8341,II27121);
  nand NAND2_5206(II27123,WX8249,II27121);
  nand NAND2_5207(WX8785,II27122,II27123);
  nand NAND2_5208(II27134,WX8342,WX8251);
  nand NAND2_5209(II27135,WX8342,II27134);
  nand NAND2_5210(II27136,WX8251,II27134);
  nand NAND2_5211(WX8792,II27135,II27136);
  nand NAND2_5212(II27147,WX8343,WX8253);
  nand NAND2_5213(II27148,WX8343,II27147);
  nand NAND2_5214(II27149,WX8253,II27147);
  nand NAND2_5215(WX8799,II27148,II27149);
  nand NAND2_5216(II27160,WX8344,WX8255);
  nand NAND2_5217(II27161,WX8344,II27160);
  nand NAND2_5218(II27162,WX8255,II27160);
  nand NAND2_5219(WX8806,II27161,II27162);
  nand NAND2_5220(II27173,WX8345,WX8257);
  nand NAND2_5221(II27174,WX8345,II27173);
  nand NAND2_5222(II27175,WX8257,II27173);
  nand NAND2_5223(WX8813,II27174,II27175);
  nand NAND2_5224(II27186,WX8346,WX8259);
  nand NAND2_5225(II27187,WX8346,II27186);
  nand NAND2_5226(II27188,WX8259,II27186);
  nand NAND2_5227(WX8820,II27187,II27188);
  nand NAND2_5228(II27199,WX8347,WX8261);
  nand NAND2_5229(II27200,WX8347,II27199);
  nand NAND2_5230(II27201,WX8261,II27199);
  nand NAND2_5231(WX8827,II27200,II27201);
  nand NAND2_5232(II27212,WX8348,WX8263);
  nand NAND2_5233(II27213,WX8348,II27212);
  nand NAND2_5234(II27214,WX8263,II27212);
  nand NAND2_5235(WX8834,II27213,II27214);
  nand NAND2_5236(II27225,WX8349,WX8265);
  nand NAND2_5237(II27226,WX8349,II27225);
  nand NAND2_5238(II27227,WX8265,II27225);
  nand NAND2_5239(WX8841,II27226,II27227);
  nand NAND2_5240(II27238,WX8350,WX8267);
  nand NAND2_5241(II27239,WX8350,II27238);
  nand NAND2_5242(II27240,WX8267,II27238);
  nand NAND2_5243(WX8848,II27239,II27240);
  nand NAND2_5244(II27251,WX8351,WX8269);
  nand NAND2_5245(II27252,WX8351,II27251);
  nand NAND2_5246(II27253,WX8269,II27251);
  nand NAND2_5247(WX8855,II27252,II27253);
  nand NAND2_5248(II27264,WX8352,WX8271);
  nand NAND2_5249(II27265,WX8352,II27264);
  nand NAND2_5250(II27266,WX8271,II27264);
  nand NAND2_5251(WX8862,II27265,II27266);
  nand NAND2_5252(II27277,WX8353,WX8273);
  nand NAND2_5253(II27278,WX8353,II27277);
  nand NAND2_5254(II27279,WX8273,II27277);
  nand NAND2_5255(WX8869,II27278,II27279);
  nand NAND2_5256(II27290,WX8354,WX8275);
  nand NAND2_5257(II27291,WX8354,II27290);
  nand NAND2_5258(II27292,WX8275,II27290);
  nand NAND2_5259(WX8876,II27291,II27292);
  nand NAND2_5260(II27303,WX8355,WX8277);
  nand NAND2_5261(II27304,WX8355,II27303);
  nand NAND2_5262(II27305,WX8277,II27303);
  nand NAND2_5263(WX8883,II27304,II27305);
  nand NAND2_5264(II27316,WX8356,WX8279);
  nand NAND2_5265(II27317,WX8356,II27316);
  nand NAND2_5266(II27318,WX8279,II27316);
  nand NAND2_5267(WX8890,II27317,II27318);
  nand NAND2_5268(II27329,WX8357,WX8281);
  nand NAND2_5269(II27330,WX8357,II27329);
  nand NAND2_5270(II27331,WX8281,II27329);
  nand NAND2_5271(WX8897,II27330,II27331);
  nand NAND2_5272(II27342,WX8358,WX8283);
  nand NAND2_5273(II27343,WX8358,II27342);
  nand NAND2_5274(II27344,WX8283,II27342);
  nand NAND2_5275(WX8904,II27343,II27344);
  nand NAND2_5276(II27355,WX8359,WX8285);
  nand NAND2_5277(II27356,WX8359,II27355);
  nand NAND2_5278(II27357,WX8285,II27355);
  nand NAND2_5279(WX8911,II27356,II27357);
  nand NAND2_5280(II27368,WX8360,WX8287);
  nand NAND2_5281(II27369,WX8360,II27368);
  nand NAND2_5282(II27370,WX8287,II27368);
  nand NAND2_5283(WX8918,II27369,II27370);
  nand NAND2_5284(II27381,WX8361,WX8289);
  nand NAND2_5285(II27382,WX8361,II27381);
  nand NAND2_5286(II27383,WX8289,II27381);
  nand NAND2_5287(WX8925,II27382,II27383);
  nand NAND2_5288(II27394,WX8362,WX8291);
  nand NAND2_5289(II27395,WX8362,II27394);
  nand NAND2_5290(II27396,WX8291,II27394);
  nand NAND2_5291(WX8932,II27395,II27396);
  nand NAND2_5292(II27407,WX8363,WX8293);
  nand NAND2_5293(II27408,WX8363,II27407);
  nand NAND2_5294(II27409,WX8293,II27407);
  nand NAND2_5295(WX8939,II27408,II27409);
  nand NAND2_5296(II27420,WX8364,WX8295);
  nand NAND2_5297(II27421,WX8364,II27420);
  nand NAND2_5298(II27422,WX8295,II27420);
  nand NAND2_5299(WX8946,II27421,II27422);
  nand NAND2_5300(II27433,WX8365,WX8297);
  nand NAND2_5301(II27434,WX8365,II27433);
  nand NAND2_5302(II27435,WX8297,II27433);
  nand NAND2_5303(WX8953,II27434,II27435);
  nand NAND2_5304(II27446,WX8366,WX8299);
  nand NAND2_5305(II27447,WX8366,II27446);
  nand NAND2_5306(II27448,WX8299,II27446);
  nand NAND2_5307(WX8960,II27447,II27448);
  nand NAND2_5308(II27459,WX8367,WX8301);
  nand NAND2_5309(II27460,WX8367,II27459);
  nand NAND2_5310(II27461,WX8301,II27459);
  nand NAND2_5311(WX8967,II27460,II27461);
  nand NAND2_5312(II27472,WX8368,WX8303);
  nand NAND2_5313(II27473,WX8368,II27472);
  nand NAND2_5314(II27474,WX8303,II27472);
  nand NAND2_5315(WX8974,II27473,II27474);
  nand NAND2_5316(II27485,WX8369,WX8305);
  nand NAND2_5317(II27486,WX8369,II27485);
  nand NAND2_5318(II27487,WX8305,II27485);
  nand NAND2_5319(WX8981,II27486,II27487);
  nand NAND2_5320(II27500,WX8385,CRC_OUT_3_31);
  nand NAND2_5321(II27501,WX8385,II27500);
  nand NAND2_5322(II27502,CRC_OUT_3_31,II27500);
  nand NAND2_5323(II27499,II27501,II27502);
  nand NAND2_5324(II27507,CRC_OUT_3_15,II27499);
  nand NAND2_5325(II27508,CRC_OUT_3_15,II27507);
  nand NAND2_5326(II27509,II27499,II27507);
  nand NAND2_5327(WX8989,II27508,II27509);
  nand NAND2_5328(II27515,WX8390,CRC_OUT_3_31);
  nand NAND2_5329(II27516,WX8390,II27515);
  nand NAND2_5330(II27517,CRC_OUT_3_31,II27515);
  nand NAND2_5331(II27514,II27516,II27517);
  nand NAND2_5332(II27522,CRC_OUT_3_10,II27514);
  nand NAND2_5333(II27523,CRC_OUT_3_10,II27522);
  nand NAND2_5334(II27524,II27514,II27522);
  nand NAND2_5335(WX8990,II27523,II27524);
  nand NAND2_5336(II27530,WX8397,CRC_OUT_3_31);
  nand NAND2_5337(II27531,WX8397,II27530);
  nand NAND2_5338(II27532,CRC_OUT_3_31,II27530);
  nand NAND2_5339(II27529,II27531,II27532);
  nand NAND2_5340(II27537,CRC_OUT_3_3,II27529);
  nand NAND2_5341(II27538,CRC_OUT_3_3,II27537);
  nand NAND2_5342(II27539,II27529,II27537);
  nand NAND2_5343(WX8991,II27538,II27539);
  nand NAND2_5344(II27544,WX8401,CRC_OUT_3_31);
  nand NAND2_5345(II27545,WX8401,II27544);
  nand NAND2_5346(II27546,CRC_OUT_3_31,II27544);
  nand NAND2_5347(WX8992,II27545,II27546);
  nand NAND2_5348(II27551,WX8370,CRC_OUT_3_30);
  nand NAND2_5349(II27552,WX8370,II27551);
  nand NAND2_5350(II27553,CRC_OUT_3_30,II27551);
  nand NAND2_5351(WX8993,II27552,II27553);
  nand NAND2_5352(II27558,WX8371,CRC_OUT_3_29);
  nand NAND2_5353(II27559,WX8371,II27558);
  nand NAND2_5354(II27560,CRC_OUT_3_29,II27558);
  nand NAND2_5355(WX8994,II27559,II27560);
  nand NAND2_5356(II27565,WX8372,CRC_OUT_3_28);
  nand NAND2_5357(II27566,WX8372,II27565);
  nand NAND2_5358(II27567,CRC_OUT_3_28,II27565);
  nand NAND2_5359(WX8995,II27566,II27567);
  nand NAND2_5360(II27572,WX8373,CRC_OUT_3_27);
  nand NAND2_5361(II27573,WX8373,II27572);
  nand NAND2_5362(II27574,CRC_OUT_3_27,II27572);
  nand NAND2_5363(WX8996,II27573,II27574);
  nand NAND2_5364(II27579,WX8374,CRC_OUT_3_26);
  nand NAND2_5365(II27580,WX8374,II27579);
  nand NAND2_5366(II27581,CRC_OUT_3_26,II27579);
  nand NAND2_5367(WX8997,II27580,II27581);
  nand NAND2_5368(II27586,WX8375,CRC_OUT_3_25);
  nand NAND2_5369(II27587,WX8375,II27586);
  nand NAND2_5370(II27588,CRC_OUT_3_25,II27586);
  nand NAND2_5371(WX8998,II27587,II27588);
  nand NAND2_5372(II27593,WX8376,CRC_OUT_3_24);
  nand NAND2_5373(II27594,WX8376,II27593);
  nand NAND2_5374(II27595,CRC_OUT_3_24,II27593);
  nand NAND2_5375(WX8999,II27594,II27595);
  nand NAND2_5376(II27600,WX8377,CRC_OUT_3_23);
  nand NAND2_5377(II27601,WX8377,II27600);
  nand NAND2_5378(II27602,CRC_OUT_3_23,II27600);
  nand NAND2_5379(WX9000,II27601,II27602);
  nand NAND2_5380(II27607,WX8378,CRC_OUT_3_22);
  nand NAND2_5381(II27608,WX8378,II27607);
  nand NAND2_5382(II27609,CRC_OUT_3_22,II27607);
  nand NAND2_5383(WX9001,II27608,II27609);
  nand NAND2_5384(II27614,WX8379,CRC_OUT_3_21);
  nand NAND2_5385(II27615,WX8379,II27614);
  nand NAND2_5386(II27616,CRC_OUT_3_21,II27614);
  nand NAND2_5387(WX9002,II27615,II27616);
  nand NAND2_5388(II27621,WX8380,CRC_OUT_3_20);
  nand NAND2_5389(II27622,WX8380,II27621);
  nand NAND2_5390(II27623,CRC_OUT_3_20,II27621);
  nand NAND2_5391(WX9003,II27622,II27623);
  nand NAND2_5392(II27628,WX8381,CRC_OUT_3_19);
  nand NAND2_5393(II27629,WX8381,II27628);
  nand NAND2_5394(II27630,CRC_OUT_3_19,II27628);
  nand NAND2_5395(WX9004,II27629,II27630);
  nand NAND2_5396(II27635,WX8382,CRC_OUT_3_18);
  nand NAND2_5397(II27636,WX8382,II27635);
  nand NAND2_5398(II27637,CRC_OUT_3_18,II27635);
  nand NAND2_5399(WX9005,II27636,II27637);
  nand NAND2_5400(II27642,WX8383,CRC_OUT_3_17);
  nand NAND2_5401(II27643,WX8383,II27642);
  nand NAND2_5402(II27644,CRC_OUT_3_17,II27642);
  nand NAND2_5403(WX9006,II27643,II27644);
  nand NAND2_5404(II27649,WX8384,CRC_OUT_3_16);
  nand NAND2_5405(II27650,WX8384,II27649);
  nand NAND2_5406(II27651,CRC_OUT_3_16,II27649);
  nand NAND2_5407(WX9007,II27650,II27651);
  nand NAND2_5408(II27656,WX8386,CRC_OUT_3_14);
  nand NAND2_5409(II27657,WX8386,II27656);
  nand NAND2_5410(II27658,CRC_OUT_3_14,II27656);
  nand NAND2_5411(WX9008,II27657,II27658);
  nand NAND2_5412(II27663,WX8387,CRC_OUT_3_13);
  nand NAND2_5413(II27664,WX8387,II27663);
  nand NAND2_5414(II27665,CRC_OUT_3_13,II27663);
  nand NAND2_5415(WX9009,II27664,II27665);
  nand NAND2_5416(II27670,WX8388,CRC_OUT_3_12);
  nand NAND2_5417(II27671,WX8388,II27670);
  nand NAND2_5418(II27672,CRC_OUT_3_12,II27670);
  nand NAND2_5419(WX9010,II27671,II27672);
  nand NAND2_5420(II27677,WX8389,CRC_OUT_3_11);
  nand NAND2_5421(II27678,WX8389,II27677);
  nand NAND2_5422(II27679,CRC_OUT_3_11,II27677);
  nand NAND2_5423(WX9011,II27678,II27679);
  nand NAND2_5424(II27684,WX8391,CRC_OUT_3_9);
  nand NAND2_5425(II27685,WX8391,II27684);
  nand NAND2_5426(II27686,CRC_OUT_3_9,II27684);
  nand NAND2_5427(WX9012,II27685,II27686);
  nand NAND2_5428(II27691,WX8392,CRC_OUT_3_8);
  nand NAND2_5429(II27692,WX8392,II27691);
  nand NAND2_5430(II27693,CRC_OUT_3_8,II27691);
  nand NAND2_5431(WX9013,II27692,II27693);
  nand NAND2_5432(II27698,WX8393,CRC_OUT_3_7);
  nand NAND2_5433(II27699,WX8393,II27698);
  nand NAND2_5434(II27700,CRC_OUT_3_7,II27698);
  nand NAND2_5435(WX9014,II27699,II27700);
  nand NAND2_5436(II27705,WX8394,CRC_OUT_3_6);
  nand NAND2_5437(II27706,WX8394,II27705);
  nand NAND2_5438(II27707,CRC_OUT_3_6,II27705);
  nand NAND2_5439(WX9015,II27706,II27707);
  nand NAND2_5440(II27712,WX8395,CRC_OUT_3_5);
  nand NAND2_5441(II27713,WX8395,II27712);
  nand NAND2_5442(II27714,CRC_OUT_3_5,II27712);
  nand NAND2_5443(WX9016,II27713,II27714);
  nand NAND2_5444(II27719,WX8396,CRC_OUT_3_4);
  nand NAND2_5445(II27720,WX8396,II27719);
  nand NAND2_5446(II27721,CRC_OUT_3_4,II27719);
  nand NAND2_5447(WX9017,II27720,II27721);
  nand NAND2_5448(II27726,WX8398,CRC_OUT_3_2);
  nand NAND2_5449(II27727,WX8398,II27726);
  nand NAND2_5450(II27728,CRC_OUT_3_2,II27726);
  nand NAND2_5451(WX9018,II27727,II27728);
  nand NAND2_5452(II27733,WX8399,CRC_OUT_3_1);
  nand NAND2_5453(II27734,WX8399,II27733);
  nand NAND2_5454(II27735,CRC_OUT_3_1,II27733);
  nand NAND2_5455(WX9019,II27734,II27735);
  nand NAND2_5456(II27740,WX8400,CRC_OUT_3_0);
  nand NAND2_5457(II27741,WX8400,II27740);
  nand NAND2_5458(II27742,CRC_OUT_3_0,II27740);
  nand NAND2_5459(WX9020,II27741,II27742);
  nand NAND2_5460(II30023,WX10052,WX9696);
  nand NAND2_5461(II30024,WX10052,II30023);
  nand NAND2_5462(II30025,WX9696,II30023);
  nand NAND2_5463(II30022,II30024,II30025);
  nand NAND2_5464(II30030,WX9760,II30022);
  nand NAND2_5465(II30031,WX9760,II30030);
  nand NAND2_5466(II30032,II30022,II30030);
  nand NAND2_5467(II30021,II30031,II30032);
  nand NAND2_5468(II30038,WX9824,WX9888);
  nand NAND2_5469(II30039,WX9824,II30038);
  nand NAND2_5470(II30040,WX9888,II30038);
  nand NAND2_5471(II30037,II30039,II30040);
  nand NAND2_5472(II30045,II30021,II30037);
  nand NAND2_5473(II30046,II30021,II30045);
  nand NAND2_5474(II30047,II30037,II30045);
  nand NAND2_5475(WX9951,II30046,II30047);
  nand NAND2_5476(II30054,WX10052,WX9698);
  nand NAND2_5477(II30055,WX10052,II30054);
  nand NAND2_5478(II30056,WX9698,II30054);
  nand NAND2_5479(II30053,II30055,II30056);
  nand NAND2_5480(II30061,WX9762,II30053);
  nand NAND2_5481(II30062,WX9762,II30061);
  nand NAND2_5482(II30063,II30053,II30061);
  nand NAND2_5483(II30052,II30062,II30063);
  nand NAND2_5484(II30069,WX9826,WX9890);
  nand NAND2_5485(II30070,WX9826,II30069);
  nand NAND2_5486(II30071,WX9890,II30069);
  nand NAND2_5487(II30068,II30070,II30071);
  nand NAND2_5488(II30076,II30052,II30068);
  nand NAND2_5489(II30077,II30052,II30076);
  nand NAND2_5490(II30078,II30068,II30076);
  nand NAND2_5491(WX9952,II30077,II30078);
  nand NAND2_5492(II30085,WX10052,WX9700);
  nand NAND2_5493(II30086,WX10052,II30085);
  nand NAND2_5494(II30087,WX9700,II30085);
  nand NAND2_5495(II30084,II30086,II30087);
  nand NAND2_5496(II30092,WX9764,II30084);
  nand NAND2_5497(II30093,WX9764,II30092);
  nand NAND2_5498(II30094,II30084,II30092);
  nand NAND2_5499(II30083,II30093,II30094);
  nand NAND2_5500(II30100,WX9828,WX9892);
  nand NAND2_5501(II30101,WX9828,II30100);
  nand NAND2_5502(II30102,WX9892,II30100);
  nand NAND2_5503(II30099,II30101,II30102);
  nand NAND2_5504(II30107,II30083,II30099);
  nand NAND2_5505(II30108,II30083,II30107);
  nand NAND2_5506(II30109,II30099,II30107);
  nand NAND2_5507(WX9953,II30108,II30109);
  nand NAND2_5508(II30116,WX10052,WX9702);
  nand NAND2_5509(II30117,WX10052,II30116);
  nand NAND2_5510(II30118,WX9702,II30116);
  nand NAND2_5511(II30115,II30117,II30118);
  nand NAND2_5512(II30123,WX9766,II30115);
  nand NAND2_5513(II30124,WX9766,II30123);
  nand NAND2_5514(II30125,II30115,II30123);
  nand NAND2_5515(II30114,II30124,II30125);
  nand NAND2_5516(II30131,WX9830,WX9894);
  nand NAND2_5517(II30132,WX9830,II30131);
  nand NAND2_5518(II30133,WX9894,II30131);
  nand NAND2_5519(II30130,II30132,II30133);
  nand NAND2_5520(II30138,II30114,II30130);
  nand NAND2_5521(II30139,II30114,II30138);
  nand NAND2_5522(II30140,II30130,II30138);
  nand NAND2_5523(WX9954,II30139,II30140);
  nand NAND2_5524(II30147,WX10052,WX9704);
  nand NAND2_5525(II30148,WX10052,II30147);
  nand NAND2_5526(II30149,WX9704,II30147);
  nand NAND2_5527(II30146,II30148,II30149);
  nand NAND2_5528(II30154,WX9768,II30146);
  nand NAND2_5529(II30155,WX9768,II30154);
  nand NAND2_5530(II30156,II30146,II30154);
  nand NAND2_5531(II30145,II30155,II30156);
  nand NAND2_5532(II30162,WX9832,WX9896);
  nand NAND2_5533(II30163,WX9832,II30162);
  nand NAND2_5534(II30164,WX9896,II30162);
  nand NAND2_5535(II30161,II30163,II30164);
  nand NAND2_5536(II30169,II30145,II30161);
  nand NAND2_5537(II30170,II30145,II30169);
  nand NAND2_5538(II30171,II30161,II30169);
  nand NAND2_5539(WX9955,II30170,II30171);
  nand NAND2_5540(II30178,WX10052,WX9706);
  nand NAND2_5541(II30179,WX10052,II30178);
  nand NAND2_5542(II30180,WX9706,II30178);
  nand NAND2_5543(II30177,II30179,II30180);
  nand NAND2_5544(II30185,WX9770,II30177);
  nand NAND2_5545(II30186,WX9770,II30185);
  nand NAND2_5546(II30187,II30177,II30185);
  nand NAND2_5547(II30176,II30186,II30187);
  nand NAND2_5548(II30193,WX9834,WX9898);
  nand NAND2_5549(II30194,WX9834,II30193);
  nand NAND2_5550(II30195,WX9898,II30193);
  nand NAND2_5551(II30192,II30194,II30195);
  nand NAND2_5552(II30200,II30176,II30192);
  nand NAND2_5553(II30201,II30176,II30200);
  nand NAND2_5554(II30202,II30192,II30200);
  nand NAND2_5555(WX9956,II30201,II30202);
  nand NAND2_5556(II30209,WX10052,WX9708);
  nand NAND2_5557(II30210,WX10052,II30209);
  nand NAND2_5558(II30211,WX9708,II30209);
  nand NAND2_5559(II30208,II30210,II30211);
  nand NAND2_5560(II30216,WX9772,II30208);
  nand NAND2_5561(II30217,WX9772,II30216);
  nand NAND2_5562(II30218,II30208,II30216);
  nand NAND2_5563(II30207,II30217,II30218);
  nand NAND2_5564(II30224,WX9836,WX9900);
  nand NAND2_5565(II30225,WX9836,II30224);
  nand NAND2_5566(II30226,WX9900,II30224);
  nand NAND2_5567(II30223,II30225,II30226);
  nand NAND2_5568(II30231,II30207,II30223);
  nand NAND2_5569(II30232,II30207,II30231);
  nand NAND2_5570(II30233,II30223,II30231);
  nand NAND2_5571(WX9957,II30232,II30233);
  nand NAND2_5572(II30240,WX10052,WX9710);
  nand NAND2_5573(II30241,WX10052,II30240);
  nand NAND2_5574(II30242,WX9710,II30240);
  nand NAND2_5575(II30239,II30241,II30242);
  nand NAND2_5576(II30247,WX9774,II30239);
  nand NAND2_5577(II30248,WX9774,II30247);
  nand NAND2_5578(II30249,II30239,II30247);
  nand NAND2_5579(II30238,II30248,II30249);
  nand NAND2_5580(II30255,WX9838,WX9902);
  nand NAND2_5581(II30256,WX9838,II30255);
  nand NAND2_5582(II30257,WX9902,II30255);
  nand NAND2_5583(II30254,II30256,II30257);
  nand NAND2_5584(II30262,II30238,II30254);
  nand NAND2_5585(II30263,II30238,II30262);
  nand NAND2_5586(II30264,II30254,II30262);
  nand NAND2_5587(WX9958,II30263,II30264);
  nand NAND2_5588(II30271,WX10052,WX9712);
  nand NAND2_5589(II30272,WX10052,II30271);
  nand NAND2_5590(II30273,WX9712,II30271);
  nand NAND2_5591(II30270,II30272,II30273);
  nand NAND2_5592(II30278,WX9776,II30270);
  nand NAND2_5593(II30279,WX9776,II30278);
  nand NAND2_5594(II30280,II30270,II30278);
  nand NAND2_5595(II30269,II30279,II30280);
  nand NAND2_5596(II30286,WX9840,WX9904);
  nand NAND2_5597(II30287,WX9840,II30286);
  nand NAND2_5598(II30288,WX9904,II30286);
  nand NAND2_5599(II30285,II30287,II30288);
  nand NAND2_5600(II30293,II30269,II30285);
  nand NAND2_5601(II30294,II30269,II30293);
  nand NAND2_5602(II30295,II30285,II30293);
  nand NAND2_5603(WX9959,II30294,II30295);
  nand NAND2_5604(II30302,WX10052,WX9714);
  nand NAND2_5605(II30303,WX10052,II30302);
  nand NAND2_5606(II30304,WX9714,II30302);
  nand NAND2_5607(II30301,II30303,II30304);
  nand NAND2_5608(II30309,WX9778,II30301);
  nand NAND2_5609(II30310,WX9778,II30309);
  nand NAND2_5610(II30311,II30301,II30309);
  nand NAND2_5611(II30300,II30310,II30311);
  nand NAND2_5612(II30317,WX9842,WX9906);
  nand NAND2_5613(II30318,WX9842,II30317);
  nand NAND2_5614(II30319,WX9906,II30317);
  nand NAND2_5615(II30316,II30318,II30319);
  nand NAND2_5616(II30324,II30300,II30316);
  nand NAND2_5617(II30325,II30300,II30324);
  nand NAND2_5618(II30326,II30316,II30324);
  nand NAND2_5619(WX9960,II30325,II30326);
  nand NAND2_5620(II30333,WX10052,WX9716);
  nand NAND2_5621(II30334,WX10052,II30333);
  nand NAND2_5622(II30335,WX9716,II30333);
  nand NAND2_5623(II30332,II30334,II30335);
  nand NAND2_5624(II30340,WX9780,II30332);
  nand NAND2_5625(II30341,WX9780,II30340);
  nand NAND2_5626(II30342,II30332,II30340);
  nand NAND2_5627(II30331,II30341,II30342);
  nand NAND2_5628(II30348,WX9844,WX9908);
  nand NAND2_5629(II30349,WX9844,II30348);
  nand NAND2_5630(II30350,WX9908,II30348);
  nand NAND2_5631(II30347,II30349,II30350);
  nand NAND2_5632(II30355,II30331,II30347);
  nand NAND2_5633(II30356,II30331,II30355);
  nand NAND2_5634(II30357,II30347,II30355);
  nand NAND2_5635(WX9961,II30356,II30357);
  nand NAND2_5636(II30364,WX10052,WX9718);
  nand NAND2_5637(II30365,WX10052,II30364);
  nand NAND2_5638(II30366,WX9718,II30364);
  nand NAND2_5639(II30363,II30365,II30366);
  nand NAND2_5640(II30371,WX9782,II30363);
  nand NAND2_5641(II30372,WX9782,II30371);
  nand NAND2_5642(II30373,II30363,II30371);
  nand NAND2_5643(II30362,II30372,II30373);
  nand NAND2_5644(II30379,WX9846,WX9910);
  nand NAND2_5645(II30380,WX9846,II30379);
  nand NAND2_5646(II30381,WX9910,II30379);
  nand NAND2_5647(II30378,II30380,II30381);
  nand NAND2_5648(II30386,II30362,II30378);
  nand NAND2_5649(II30387,II30362,II30386);
  nand NAND2_5650(II30388,II30378,II30386);
  nand NAND2_5651(WX9962,II30387,II30388);
  nand NAND2_5652(II30395,WX10052,WX9720);
  nand NAND2_5653(II30396,WX10052,II30395);
  nand NAND2_5654(II30397,WX9720,II30395);
  nand NAND2_5655(II30394,II30396,II30397);
  nand NAND2_5656(II30402,WX9784,II30394);
  nand NAND2_5657(II30403,WX9784,II30402);
  nand NAND2_5658(II30404,II30394,II30402);
  nand NAND2_5659(II30393,II30403,II30404);
  nand NAND2_5660(II30410,WX9848,WX9912);
  nand NAND2_5661(II30411,WX9848,II30410);
  nand NAND2_5662(II30412,WX9912,II30410);
  nand NAND2_5663(II30409,II30411,II30412);
  nand NAND2_5664(II30417,II30393,II30409);
  nand NAND2_5665(II30418,II30393,II30417);
  nand NAND2_5666(II30419,II30409,II30417);
  nand NAND2_5667(WX9963,II30418,II30419);
  nand NAND2_5668(II30426,WX10052,WX9722);
  nand NAND2_5669(II30427,WX10052,II30426);
  nand NAND2_5670(II30428,WX9722,II30426);
  nand NAND2_5671(II30425,II30427,II30428);
  nand NAND2_5672(II30433,WX9786,II30425);
  nand NAND2_5673(II30434,WX9786,II30433);
  nand NAND2_5674(II30435,II30425,II30433);
  nand NAND2_5675(II30424,II30434,II30435);
  nand NAND2_5676(II30441,WX9850,WX9914);
  nand NAND2_5677(II30442,WX9850,II30441);
  nand NAND2_5678(II30443,WX9914,II30441);
  nand NAND2_5679(II30440,II30442,II30443);
  nand NAND2_5680(II30448,II30424,II30440);
  nand NAND2_5681(II30449,II30424,II30448);
  nand NAND2_5682(II30450,II30440,II30448);
  nand NAND2_5683(WX9964,II30449,II30450);
  nand NAND2_5684(II30457,WX10052,WX9724);
  nand NAND2_5685(II30458,WX10052,II30457);
  nand NAND2_5686(II30459,WX9724,II30457);
  nand NAND2_5687(II30456,II30458,II30459);
  nand NAND2_5688(II30464,WX9788,II30456);
  nand NAND2_5689(II30465,WX9788,II30464);
  nand NAND2_5690(II30466,II30456,II30464);
  nand NAND2_5691(II30455,II30465,II30466);
  nand NAND2_5692(II30472,WX9852,WX9916);
  nand NAND2_5693(II30473,WX9852,II30472);
  nand NAND2_5694(II30474,WX9916,II30472);
  nand NAND2_5695(II30471,II30473,II30474);
  nand NAND2_5696(II30479,II30455,II30471);
  nand NAND2_5697(II30480,II30455,II30479);
  nand NAND2_5698(II30481,II30471,II30479);
  nand NAND2_5699(WX9965,II30480,II30481);
  nand NAND2_5700(II30488,WX10052,WX9726);
  nand NAND2_5701(II30489,WX10052,II30488);
  nand NAND2_5702(II30490,WX9726,II30488);
  nand NAND2_5703(II30487,II30489,II30490);
  nand NAND2_5704(II30495,WX9790,II30487);
  nand NAND2_5705(II30496,WX9790,II30495);
  nand NAND2_5706(II30497,II30487,II30495);
  nand NAND2_5707(II30486,II30496,II30497);
  nand NAND2_5708(II30503,WX9854,WX9918);
  nand NAND2_5709(II30504,WX9854,II30503);
  nand NAND2_5710(II30505,WX9918,II30503);
  nand NAND2_5711(II30502,II30504,II30505);
  nand NAND2_5712(II30510,II30486,II30502);
  nand NAND2_5713(II30511,II30486,II30510);
  nand NAND2_5714(II30512,II30502,II30510);
  nand NAND2_5715(WX9966,II30511,II30512);
  nand NAND2_5716(II30519,WX10053,WX9728);
  nand NAND2_5717(II30520,WX10053,II30519);
  nand NAND2_5718(II30521,WX9728,II30519);
  nand NAND2_5719(II30518,II30520,II30521);
  nand NAND2_5720(II30526,WX9792,II30518);
  nand NAND2_5721(II30527,WX9792,II30526);
  nand NAND2_5722(II30528,II30518,II30526);
  nand NAND2_5723(II30517,II30527,II30528);
  nand NAND2_5724(II30534,WX9856,WX9920);
  nand NAND2_5725(II30535,WX9856,II30534);
  nand NAND2_5726(II30536,WX9920,II30534);
  nand NAND2_5727(II30533,II30535,II30536);
  nand NAND2_5728(II30541,II30517,II30533);
  nand NAND2_5729(II30542,II30517,II30541);
  nand NAND2_5730(II30543,II30533,II30541);
  nand NAND2_5731(WX9967,II30542,II30543);
  nand NAND2_5732(II30550,WX10053,WX9730);
  nand NAND2_5733(II30551,WX10053,II30550);
  nand NAND2_5734(II30552,WX9730,II30550);
  nand NAND2_5735(II30549,II30551,II30552);
  nand NAND2_5736(II30557,WX9794,II30549);
  nand NAND2_5737(II30558,WX9794,II30557);
  nand NAND2_5738(II30559,II30549,II30557);
  nand NAND2_5739(II30548,II30558,II30559);
  nand NAND2_5740(II30565,WX9858,WX9922);
  nand NAND2_5741(II30566,WX9858,II30565);
  nand NAND2_5742(II30567,WX9922,II30565);
  nand NAND2_5743(II30564,II30566,II30567);
  nand NAND2_5744(II30572,II30548,II30564);
  nand NAND2_5745(II30573,II30548,II30572);
  nand NAND2_5746(II30574,II30564,II30572);
  nand NAND2_5747(WX9968,II30573,II30574);
  nand NAND2_5748(II30581,WX10053,WX9732);
  nand NAND2_5749(II30582,WX10053,II30581);
  nand NAND2_5750(II30583,WX9732,II30581);
  nand NAND2_5751(II30580,II30582,II30583);
  nand NAND2_5752(II30588,WX9796,II30580);
  nand NAND2_5753(II30589,WX9796,II30588);
  nand NAND2_5754(II30590,II30580,II30588);
  nand NAND2_5755(II30579,II30589,II30590);
  nand NAND2_5756(II30596,WX9860,WX9924);
  nand NAND2_5757(II30597,WX9860,II30596);
  nand NAND2_5758(II30598,WX9924,II30596);
  nand NAND2_5759(II30595,II30597,II30598);
  nand NAND2_5760(II30603,II30579,II30595);
  nand NAND2_5761(II30604,II30579,II30603);
  nand NAND2_5762(II30605,II30595,II30603);
  nand NAND2_5763(WX9969,II30604,II30605);
  nand NAND2_5764(II30612,WX10053,WX9734);
  nand NAND2_5765(II30613,WX10053,II30612);
  nand NAND2_5766(II30614,WX9734,II30612);
  nand NAND2_5767(II30611,II30613,II30614);
  nand NAND2_5768(II30619,WX9798,II30611);
  nand NAND2_5769(II30620,WX9798,II30619);
  nand NAND2_5770(II30621,II30611,II30619);
  nand NAND2_5771(II30610,II30620,II30621);
  nand NAND2_5772(II30627,WX9862,WX9926);
  nand NAND2_5773(II30628,WX9862,II30627);
  nand NAND2_5774(II30629,WX9926,II30627);
  nand NAND2_5775(II30626,II30628,II30629);
  nand NAND2_5776(II30634,II30610,II30626);
  nand NAND2_5777(II30635,II30610,II30634);
  nand NAND2_5778(II30636,II30626,II30634);
  nand NAND2_5779(WX9970,II30635,II30636);
  nand NAND2_5780(II30643,WX10053,WX9736);
  nand NAND2_5781(II30644,WX10053,II30643);
  nand NAND2_5782(II30645,WX9736,II30643);
  nand NAND2_5783(II30642,II30644,II30645);
  nand NAND2_5784(II30650,WX9800,II30642);
  nand NAND2_5785(II30651,WX9800,II30650);
  nand NAND2_5786(II30652,II30642,II30650);
  nand NAND2_5787(II30641,II30651,II30652);
  nand NAND2_5788(II30658,WX9864,WX9928);
  nand NAND2_5789(II30659,WX9864,II30658);
  nand NAND2_5790(II30660,WX9928,II30658);
  nand NAND2_5791(II30657,II30659,II30660);
  nand NAND2_5792(II30665,II30641,II30657);
  nand NAND2_5793(II30666,II30641,II30665);
  nand NAND2_5794(II30667,II30657,II30665);
  nand NAND2_5795(WX9971,II30666,II30667);
  nand NAND2_5796(II30674,WX10053,WX9738);
  nand NAND2_5797(II30675,WX10053,II30674);
  nand NAND2_5798(II30676,WX9738,II30674);
  nand NAND2_5799(II30673,II30675,II30676);
  nand NAND2_5800(II30681,WX9802,II30673);
  nand NAND2_5801(II30682,WX9802,II30681);
  nand NAND2_5802(II30683,II30673,II30681);
  nand NAND2_5803(II30672,II30682,II30683);
  nand NAND2_5804(II30689,WX9866,WX9930);
  nand NAND2_5805(II30690,WX9866,II30689);
  nand NAND2_5806(II30691,WX9930,II30689);
  nand NAND2_5807(II30688,II30690,II30691);
  nand NAND2_5808(II30696,II30672,II30688);
  nand NAND2_5809(II30697,II30672,II30696);
  nand NAND2_5810(II30698,II30688,II30696);
  nand NAND2_5811(WX9972,II30697,II30698);
  nand NAND2_5812(II30705,WX10053,WX9740);
  nand NAND2_5813(II30706,WX10053,II30705);
  nand NAND2_5814(II30707,WX9740,II30705);
  nand NAND2_5815(II30704,II30706,II30707);
  nand NAND2_5816(II30712,WX9804,II30704);
  nand NAND2_5817(II30713,WX9804,II30712);
  nand NAND2_5818(II30714,II30704,II30712);
  nand NAND2_5819(II30703,II30713,II30714);
  nand NAND2_5820(II30720,WX9868,WX9932);
  nand NAND2_5821(II30721,WX9868,II30720);
  nand NAND2_5822(II30722,WX9932,II30720);
  nand NAND2_5823(II30719,II30721,II30722);
  nand NAND2_5824(II30727,II30703,II30719);
  nand NAND2_5825(II30728,II30703,II30727);
  nand NAND2_5826(II30729,II30719,II30727);
  nand NAND2_5827(WX9973,II30728,II30729);
  nand NAND2_5828(II30736,WX10053,WX9742);
  nand NAND2_5829(II30737,WX10053,II30736);
  nand NAND2_5830(II30738,WX9742,II30736);
  nand NAND2_5831(II30735,II30737,II30738);
  nand NAND2_5832(II30743,WX9806,II30735);
  nand NAND2_5833(II30744,WX9806,II30743);
  nand NAND2_5834(II30745,II30735,II30743);
  nand NAND2_5835(II30734,II30744,II30745);
  nand NAND2_5836(II30751,WX9870,WX9934);
  nand NAND2_5837(II30752,WX9870,II30751);
  nand NAND2_5838(II30753,WX9934,II30751);
  nand NAND2_5839(II30750,II30752,II30753);
  nand NAND2_5840(II30758,II30734,II30750);
  nand NAND2_5841(II30759,II30734,II30758);
  nand NAND2_5842(II30760,II30750,II30758);
  nand NAND2_5843(WX9974,II30759,II30760);
  nand NAND2_5844(II30767,WX10053,WX9744);
  nand NAND2_5845(II30768,WX10053,II30767);
  nand NAND2_5846(II30769,WX9744,II30767);
  nand NAND2_5847(II30766,II30768,II30769);
  nand NAND2_5848(II30774,WX9808,II30766);
  nand NAND2_5849(II30775,WX9808,II30774);
  nand NAND2_5850(II30776,II30766,II30774);
  nand NAND2_5851(II30765,II30775,II30776);
  nand NAND2_5852(II30782,WX9872,WX9936);
  nand NAND2_5853(II30783,WX9872,II30782);
  nand NAND2_5854(II30784,WX9936,II30782);
  nand NAND2_5855(II30781,II30783,II30784);
  nand NAND2_5856(II30789,II30765,II30781);
  nand NAND2_5857(II30790,II30765,II30789);
  nand NAND2_5858(II30791,II30781,II30789);
  nand NAND2_5859(WX9975,II30790,II30791);
  nand NAND2_5860(II30798,WX10053,WX9746);
  nand NAND2_5861(II30799,WX10053,II30798);
  nand NAND2_5862(II30800,WX9746,II30798);
  nand NAND2_5863(II30797,II30799,II30800);
  nand NAND2_5864(II30805,WX9810,II30797);
  nand NAND2_5865(II30806,WX9810,II30805);
  nand NAND2_5866(II30807,II30797,II30805);
  nand NAND2_5867(II30796,II30806,II30807);
  nand NAND2_5868(II30813,WX9874,WX9938);
  nand NAND2_5869(II30814,WX9874,II30813);
  nand NAND2_5870(II30815,WX9938,II30813);
  nand NAND2_5871(II30812,II30814,II30815);
  nand NAND2_5872(II30820,II30796,II30812);
  nand NAND2_5873(II30821,II30796,II30820);
  nand NAND2_5874(II30822,II30812,II30820);
  nand NAND2_5875(WX9976,II30821,II30822);
  nand NAND2_5876(II30829,WX10053,WX9748);
  nand NAND2_5877(II30830,WX10053,II30829);
  nand NAND2_5878(II30831,WX9748,II30829);
  nand NAND2_5879(II30828,II30830,II30831);
  nand NAND2_5880(II30836,WX9812,II30828);
  nand NAND2_5881(II30837,WX9812,II30836);
  nand NAND2_5882(II30838,II30828,II30836);
  nand NAND2_5883(II30827,II30837,II30838);
  nand NAND2_5884(II30844,WX9876,WX9940);
  nand NAND2_5885(II30845,WX9876,II30844);
  nand NAND2_5886(II30846,WX9940,II30844);
  nand NAND2_5887(II30843,II30845,II30846);
  nand NAND2_5888(II30851,II30827,II30843);
  nand NAND2_5889(II30852,II30827,II30851);
  nand NAND2_5890(II30853,II30843,II30851);
  nand NAND2_5891(WX9977,II30852,II30853);
  nand NAND2_5892(II30860,WX10053,WX9750);
  nand NAND2_5893(II30861,WX10053,II30860);
  nand NAND2_5894(II30862,WX9750,II30860);
  nand NAND2_5895(II30859,II30861,II30862);
  nand NAND2_5896(II30867,WX9814,II30859);
  nand NAND2_5897(II30868,WX9814,II30867);
  nand NAND2_5898(II30869,II30859,II30867);
  nand NAND2_5899(II30858,II30868,II30869);
  nand NAND2_5900(II30875,WX9878,WX9942);
  nand NAND2_5901(II30876,WX9878,II30875);
  nand NAND2_5902(II30877,WX9942,II30875);
  nand NAND2_5903(II30874,II30876,II30877);
  nand NAND2_5904(II30882,II30858,II30874);
  nand NAND2_5905(II30883,II30858,II30882);
  nand NAND2_5906(II30884,II30874,II30882);
  nand NAND2_5907(WX9978,II30883,II30884);
  nand NAND2_5908(II30891,WX10053,WX9752);
  nand NAND2_5909(II30892,WX10053,II30891);
  nand NAND2_5910(II30893,WX9752,II30891);
  nand NAND2_5911(II30890,II30892,II30893);
  nand NAND2_5912(II30898,WX9816,II30890);
  nand NAND2_5913(II30899,WX9816,II30898);
  nand NAND2_5914(II30900,II30890,II30898);
  nand NAND2_5915(II30889,II30899,II30900);
  nand NAND2_5916(II30906,WX9880,WX9944);
  nand NAND2_5917(II30907,WX9880,II30906);
  nand NAND2_5918(II30908,WX9944,II30906);
  nand NAND2_5919(II30905,II30907,II30908);
  nand NAND2_5920(II30913,II30889,II30905);
  nand NAND2_5921(II30914,II30889,II30913);
  nand NAND2_5922(II30915,II30905,II30913);
  nand NAND2_5923(WX9979,II30914,II30915);
  nand NAND2_5924(II30922,WX10053,WX9754);
  nand NAND2_5925(II30923,WX10053,II30922);
  nand NAND2_5926(II30924,WX9754,II30922);
  nand NAND2_5927(II30921,II30923,II30924);
  nand NAND2_5928(II30929,WX9818,II30921);
  nand NAND2_5929(II30930,WX9818,II30929);
  nand NAND2_5930(II30931,II30921,II30929);
  nand NAND2_5931(II30920,II30930,II30931);
  nand NAND2_5932(II30937,WX9882,WX9946);
  nand NAND2_5933(II30938,WX9882,II30937);
  nand NAND2_5934(II30939,WX9946,II30937);
  nand NAND2_5935(II30936,II30938,II30939);
  nand NAND2_5936(II30944,II30920,II30936);
  nand NAND2_5937(II30945,II30920,II30944);
  nand NAND2_5938(II30946,II30936,II30944);
  nand NAND2_5939(WX9980,II30945,II30946);
  nand NAND2_5940(II30953,WX10053,WX9756);
  nand NAND2_5941(II30954,WX10053,II30953);
  nand NAND2_5942(II30955,WX9756,II30953);
  nand NAND2_5943(II30952,II30954,II30955);
  nand NAND2_5944(II30960,WX9820,II30952);
  nand NAND2_5945(II30961,WX9820,II30960);
  nand NAND2_5946(II30962,II30952,II30960);
  nand NAND2_5947(II30951,II30961,II30962);
  nand NAND2_5948(II30968,WX9884,WX9948);
  nand NAND2_5949(II30969,WX9884,II30968);
  nand NAND2_5950(II30970,WX9948,II30968);
  nand NAND2_5951(II30967,II30969,II30970);
  nand NAND2_5952(II30975,II30951,II30967);
  nand NAND2_5953(II30976,II30951,II30975);
  nand NAND2_5954(II30977,II30967,II30975);
  nand NAND2_5955(WX9981,II30976,II30977);
  nand NAND2_5956(II30984,WX10053,WX9758);
  nand NAND2_5957(II30985,WX10053,II30984);
  nand NAND2_5958(II30986,WX9758,II30984);
  nand NAND2_5959(II30983,II30985,II30986);
  nand NAND2_5960(II30991,WX9822,II30983);
  nand NAND2_5961(II30992,WX9822,II30991);
  nand NAND2_5962(II30993,II30983,II30991);
  nand NAND2_5963(II30982,II30992,II30993);
  nand NAND2_5964(II30999,WX9886,WX9950);
  nand NAND2_5965(II31000,WX9886,II30999);
  nand NAND2_5966(II31001,WX9950,II30999);
  nand NAND2_5967(II30998,II31000,II31001);
  nand NAND2_5968(II31006,II30982,II30998);
  nand NAND2_5969(II31007,II30982,II31006);
  nand NAND2_5970(II31008,II30998,II31006);
  nand NAND2_5971(WX9982,II31007,II31008);
  nand NAND2_5972(II31087,WX9631,WX9536);
  nand NAND2_5973(II31088,WX9631,II31087);
  nand NAND2_5974(II31089,WX9536,II31087);
  nand NAND2_5975(WX10057,II31088,II31089);
  nand NAND2_5976(II31100,WX9632,WX9538);
  nand NAND2_5977(II31101,WX9632,II31100);
  nand NAND2_5978(II31102,WX9538,II31100);
  nand NAND2_5979(WX10064,II31101,II31102);
  nand NAND2_5980(II31113,WX9633,WX9540);
  nand NAND2_5981(II31114,WX9633,II31113);
  nand NAND2_5982(II31115,WX9540,II31113);
  nand NAND2_5983(WX10071,II31114,II31115);
  nand NAND2_5984(II31126,WX9634,WX9542);
  nand NAND2_5985(II31127,WX9634,II31126);
  nand NAND2_5986(II31128,WX9542,II31126);
  nand NAND2_5987(WX10078,II31127,II31128);
  nand NAND2_5988(II31139,WX9635,WX9544);
  nand NAND2_5989(II31140,WX9635,II31139);
  nand NAND2_5990(II31141,WX9544,II31139);
  nand NAND2_5991(WX10085,II31140,II31141);
  nand NAND2_5992(II31152,WX9636,WX9546);
  nand NAND2_5993(II31153,WX9636,II31152);
  nand NAND2_5994(II31154,WX9546,II31152);
  nand NAND2_5995(WX10092,II31153,II31154);
  nand NAND2_5996(II31165,WX9637,WX9548);
  nand NAND2_5997(II31166,WX9637,II31165);
  nand NAND2_5998(II31167,WX9548,II31165);
  nand NAND2_5999(WX10099,II31166,II31167);
  nand NAND2_6000(II31178,WX9638,WX9550);
  nand NAND2_6001(II31179,WX9638,II31178);
  nand NAND2_6002(II31180,WX9550,II31178);
  nand NAND2_6003(WX10106,II31179,II31180);
  nand NAND2_6004(II31191,WX9639,WX9552);
  nand NAND2_6005(II31192,WX9639,II31191);
  nand NAND2_6006(II31193,WX9552,II31191);
  nand NAND2_6007(WX10113,II31192,II31193);
  nand NAND2_6008(II31204,WX9640,WX9554);
  nand NAND2_6009(II31205,WX9640,II31204);
  nand NAND2_6010(II31206,WX9554,II31204);
  nand NAND2_6011(WX10120,II31205,II31206);
  nand NAND2_6012(II31217,WX9641,WX9556);
  nand NAND2_6013(II31218,WX9641,II31217);
  nand NAND2_6014(II31219,WX9556,II31217);
  nand NAND2_6015(WX10127,II31218,II31219);
  nand NAND2_6016(II31230,WX9642,WX9558);
  nand NAND2_6017(II31231,WX9642,II31230);
  nand NAND2_6018(II31232,WX9558,II31230);
  nand NAND2_6019(WX10134,II31231,II31232);
  nand NAND2_6020(II31243,WX9643,WX9560);
  nand NAND2_6021(II31244,WX9643,II31243);
  nand NAND2_6022(II31245,WX9560,II31243);
  nand NAND2_6023(WX10141,II31244,II31245);
  nand NAND2_6024(II31256,WX9644,WX9562);
  nand NAND2_6025(II31257,WX9644,II31256);
  nand NAND2_6026(II31258,WX9562,II31256);
  nand NAND2_6027(WX10148,II31257,II31258);
  nand NAND2_6028(II31269,WX9645,WX9564);
  nand NAND2_6029(II31270,WX9645,II31269);
  nand NAND2_6030(II31271,WX9564,II31269);
  nand NAND2_6031(WX10155,II31270,II31271);
  nand NAND2_6032(II31282,WX9646,WX9566);
  nand NAND2_6033(II31283,WX9646,II31282);
  nand NAND2_6034(II31284,WX9566,II31282);
  nand NAND2_6035(WX10162,II31283,II31284);
  nand NAND2_6036(II31295,WX9647,WX9568);
  nand NAND2_6037(II31296,WX9647,II31295);
  nand NAND2_6038(II31297,WX9568,II31295);
  nand NAND2_6039(WX10169,II31296,II31297);
  nand NAND2_6040(II31308,WX9648,WX9570);
  nand NAND2_6041(II31309,WX9648,II31308);
  nand NAND2_6042(II31310,WX9570,II31308);
  nand NAND2_6043(WX10176,II31309,II31310);
  nand NAND2_6044(II31321,WX9649,WX9572);
  nand NAND2_6045(II31322,WX9649,II31321);
  nand NAND2_6046(II31323,WX9572,II31321);
  nand NAND2_6047(WX10183,II31322,II31323);
  nand NAND2_6048(II31334,WX9650,WX9574);
  nand NAND2_6049(II31335,WX9650,II31334);
  nand NAND2_6050(II31336,WX9574,II31334);
  nand NAND2_6051(WX10190,II31335,II31336);
  nand NAND2_6052(II31347,WX9651,WX9576);
  nand NAND2_6053(II31348,WX9651,II31347);
  nand NAND2_6054(II31349,WX9576,II31347);
  nand NAND2_6055(WX10197,II31348,II31349);
  nand NAND2_6056(II31360,WX9652,WX9578);
  nand NAND2_6057(II31361,WX9652,II31360);
  nand NAND2_6058(II31362,WX9578,II31360);
  nand NAND2_6059(WX10204,II31361,II31362);
  nand NAND2_6060(II31373,WX9653,WX9580);
  nand NAND2_6061(II31374,WX9653,II31373);
  nand NAND2_6062(II31375,WX9580,II31373);
  nand NAND2_6063(WX10211,II31374,II31375);
  nand NAND2_6064(II31386,WX9654,WX9582);
  nand NAND2_6065(II31387,WX9654,II31386);
  nand NAND2_6066(II31388,WX9582,II31386);
  nand NAND2_6067(WX10218,II31387,II31388);
  nand NAND2_6068(II31399,WX9655,WX9584);
  nand NAND2_6069(II31400,WX9655,II31399);
  nand NAND2_6070(II31401,WX9584,II31399);
  nand NAND2_6071(WX10225,II31400,II31401);
  nand NAND2_6072(II31412,WX9656,WX9586);
  nand NAND2_6073(II31413,WX9656,II31412);
  nand NAND2_6074(II31414,WX9586,II31412);
  nand NAND2_6075(WX10232,II31413,II31414);
  nand NAND2_6076(II31425,WX9657,WX9588);
  nand NAND2_6077(II31426,WX9657,II31425);
  nand NAND2_6078(II31427,WX9588,II31425);
  nand NAND2_6079(WX10239,II31426,II31427);
  nand NAND2_6080(II31438,WX9658,WX9590);
  nand NAND2_6081(II31439,WX9658,II31438);
  nand NAND2_6082(II31440,WX9590,II31438);
  nand NAND2_6083(WX10246,II31439,II31440);
  nand NAND2_6084(II31451,WX9659,WX9592);
  nand NAND2_6085(II31452,WX9659,II31451);
  nand NAND2_6086(II31453,WX9592,II31451);
  nand NAND2_6087(WX10253,II31452,II31453);
  nand NAND2_6088(II31464,WX9660,WX9594);
  nand NAND2_6089(II31465,WX9660,II31464);
  nand NAND2_6090(II31466,WX9594,II31464);
  nand NAND2_6091(WX10260,II31465,II31466);
  nand NAND2_6092(II31477,WX9661,WX9596);
  nand NAND2_6093(II31478,WX9661,II31477);
  nand NAND2_6094(II31479,WX9596,II31477);
  nand NAND2_6095(WX10267,II31478,II31479);
  nand NAND2_6096(II31490,WX9662,WX9598);
  nand NAND2_6097(II31491,WX9662,II31490);
  nand NAND2_6098(II31492,WX9598,II31490);
  nand NAND2_6099(WX10274,II31491,II31492);
  nand NAND2_6100(II31505,WX9678,CRC_OUT_2_31);
  nand NAND2_6101(II31506,WX9678,II31505);
  nand NAND2_6102(II31507,CRC_OUT_2_31,II31505);
  nand NAND2_6103(II31504,II31506,II31507);
  nand NAND2_6104(II31512,CRC_OUT_2_15,II31504);
  nand NAND2_6105(II31513,CRC_OUT_2_15,II31512);
  nand NAND2_6106(II31514,II31504,II31512);
  nand NAND2_6107(WX10282,II31513,II31514);
  nand NAND2_6108(II31520,WX9683,CRC_OUT_2_31);
  nand NAND2_6109(II31521,WX9683,II31520);
  nand NAND2_6110(II31522,CRC_OUT_2_31,II31520);
  nand NAND2_6111(II31519,II31521,II31522);
  nand NAND2_6112(II31527,CRC_OUT_2_10,II31519);
  nand NAND2_6113(II31528,CRC_OUT_2_10,II31527);
  nand NAND2_6114(II31529,II31519,II31527);
  nand NAND2_6115(WX10283,II31528,II31529);
  nand NAND2_6116(II31535,WX9690,CRC_OUT_2_31);
  nand NAND2_6117(II31536,WX9690,II31535);
  nand NAND2_6118(II31537,CRC_OUT_2_31,II31535);
  nand NAND2_6119(II31534,II31536,II31537);
  nand NAND2_6120(II31542,CRC_OUT_2_3,II31534);
  nand NAND2_6121(II31543,CRC_OUT_2_3,II31542);
  nand NAND2_6122(II31544,II31534,II31542);
  nand NAND2_6123(WX10284,II31543,II31544);
  nand NAND2_6124(II31549,WX9694,CRC_OUT_2_31);
  nand NAND2_6125(II31550,WX9694,II31549);
  nand NAND2_6126(II31551,CRC_OUT_2_31,II31549);
  nand NAND2_6127(WX10285,II31550,II31551);
  nand NAND2_6128(II31556,WX9663,CRC_OUT_2_30);
  nand NAND2_6129(II31557,WX9663,II31556);
  nand NAND2_6130(II31558,CRC_OUT_2_30,II31556);
  nand NAND2_6131(WX10286,II31557,II31558);
  nand NAND2_6132(II31563,WX9664,CRC_OUT_2_29);
  nand NAND2_6133(II31564,WX9664,II31563);
  nand NAND2_6134(II31565,CRC_OUT_2_29,II31563);
  nand NAND2_6135(WX10287,II31564,II31565);
  nand NAND2_6136(II31570,WX9665,CRC_OUT_2_28);
  nand NAND2_6137(II31571,WX9665,II31570);
  nand NAND2_6138(II31572,CRC_OUT_2_28,II31570);
  nand NAND2_6139(WX10288,II31571,II31572);
  nand NAND2_6140(II31577,WX9666,CRC_OUT_2_27);
  nand NAND2_6141(II31578,WX9666,II31577);
  nand NAND2_6142(II31579,CRC_OUT_2_27,II31577);
  nand NAND2_6143(WX10289,II31578,II31579);
  nand NAND2_6144(II31584,WX9667,CRC_OUT_2_26);
  nand NAND2_6145(II31585,WX9667,II31584);
  nand NAND2_6146(II31586,CRC_OUT_2_26,II31584);
  nand NAND2_6147(WX10290,II31585,II31586);
  nand NAND2_6148(II31591,WX9668,CRC_OUT_2_25);
  nand NAND2_6149(II31592,WX9668,II31591);
  nand NAND2_6150(II31593,CRC_OUT_2_25,II31591);
  nand NAND2_6151(WX10291,II31592,II31593);
  nand NAND2_6152(II31598,WX9669,CRC_OUT_2_24);
  nand NAND2_6153(II31599,WX9669,II31598);
  nand NAND2_6154(II31600,CRC_OUT_2_24,II31598);
  nand NAND2_6155(WX10292,II31599,II31600);
  nand NAND2_6156(II31605,WX9670,CRC_OUT_2_23);
  nand NAND2_6157(II31606,WX9670,II31605);
  nand NAND2_6158(II31607,CRC_OUT_2_23,II31605);
  nand NAND2_6159(WX10293,II31606,II31607);
  nand NAND2_6160(II31612,WX9671,CRC_OUT_2_22);
  nand NAND2_6161(II31613,WX9671,II31612);
  nand NAND2_6162(II31614,CRC_OUT_2_22,II31612);
  nand NAND2_6163(WX10294,II31613,II31614);
  nand NAND2_6164(II31619,WX9672,CRC_OUT_2_21);
  nand NAND2_6165(II31620,WX9672,II31619);
  nand NAND2_6166(II31621,CRC_OUT_2_21,II31619);
  nand NAND2_6167(WX10295,II31620,II31621);
  nand NAND2_6168(II31626,WX9673,CRC_OUT_2_20);
  nand NAND2_6169(II31627,WX9673,II31626);
  nand NAND2_6170(II31628,CRC_OUT_2_20,II31626);
  nand NAND2_6171(WX10296,II31627,II31628);
  nand NAND2_6172(II31633,WX9674,CRC_OUT_2_19);
  nand NAND2_6173(II31634,WX9674,II31633);
  nand NAND2_6174(II31635,CRC_OUT_2_19,II31633);
  nand NAND2_6175(WX10297,II31634,II31635);
  nand NAND2_6176(II31640,WX9675,CRC_OUT_2_18);
  nand NAND2_6177(II31641,WX9675,II31640);
  nand NAND2_6178(II31642,CRC_OUT_2_18,II31640);
  nand NAND2_6179(WX10298,II31641,II31642);
  nand NAND2_6180(II31647,WX9676,CRC_OUT_2_17);
  nand NAND2_6181(II31648,WX9676,II31647);
  nand NAND2_6182(II31649,CRC_OUT_2_17,II31647);
  nand NAND2_6183(WX10299,II31648,II31649);
  nand NAND2_6184(II31654,WX9677,CRC_OUT_2_16);
  nand NAND2_6185(II31655,WX9677,II31654);
  nand NAND2_6186(II31656,CRC_OUT_2_16,II31654);
  nand NAND2_6187(WX10300,II31655,II31656);
  nand NAND2_6188(II31661,WX9679,CRC_OUT_2_14);
  nand NAND2_6189(II31662,WX9679,II31661);
  nand NAND2_6190(II31663,CRC_OUT_2_14,II31661);
  nand NAND2_6191(WX10301,II31662,II31663);
  nand NAND2_6192(II31668,WX9680,CRC_OUT_2_13);
  nand NAND2_6193(II31669,WX9680,II31668);
  nand NAND2_6194(II31670,CRC_OUT_2_13,II31668);
  nand NAND2_6195(WX10302,II31669,II31670);
  nand NAND2_6196(II31675,WX9681,CRC_OUT_2_12);
  nand NAND2_6197(II31676,WX9681,II31675);
  nand NAND2_6198(II31677,CRC_OUT_2_12,II31675);
  nand NAND2_6199(WX10303,II31676,II31677);
  nand NAND2_6200(II31682,WX9682,CRC_OUT_2_11);
  nand NAND2_6201(II31683,WX9682,II31682);
  nand NAND2_6202(II31684,CRC_OUT_2_11,II31682);
  nand NAND2_6203(WX10304,II31683,II31684);
  nand NAND2_6204(II31689,WX9684,CRC_OUT_2_9);
  nand NAND2_6205(II31690,WX9684,II31689);
  nand NAND2_6206(II31691,CRC_OUT_2_9,II31689);
  nand NAND2_6207(WX10305,II31690,II31691);
  nand NAND2_6208(II31696,WX9685,CRC_OUT_2_8);
  nand NAND2_6209(II31697,WX9685,II31696);
  nand NAND2_6210(II31698,CRC_OUT_2_8,II31696);
  nand NAND2_6211(WX10306,II31697,II31698);
  nand NAND2_6212(II31703,WX9686,CRC_OUT_2_7);
  nand NAND2_6213(II31704,WX9686,II31703);
  nand NAND2_6214(II31705,CRC_OUT_2_7,II31703);
  nand NAND2_6215(WX10307,II31704,II31705);
  nand NAND2_6216(II31710,WX9687,CRC_OUT_2_6);
  nand NAND2_6217(II31711,WX9687,II31710);
  nand NAND2_6218(II31712,CRC_OUT_2_6,II31710);
  nand NAND2_6219(WX10308,II31711,II31712);
  nand NAND2_6220(II31717,WX9688,CRC_OUT_2_5);
  nand NAND2_6221(II31718,WX9688,II31717);
  nand NAND2_6222(II31719,CRC_OUT_2_5,II31717);
  nand NAND2_6223(WX10309,II31718,II31719);
  nand NAND2_6224(II31724,WX9689,CRC_OUT_2_4);
  nand NAND2_6225(II31725,WX9689,II31724);
  nand NAND2_6226(II31726,CRC_OUT_2_4,II31724);
  nand NAND2_6227(WX10310,II31725,II31726);
  nand NAND2_6228(II31731,WX9691,CRC_OUT_2_2);
  nand NAND2_6229(II31732,WX9691,II31731);
  nand NAND2_6230(II31733,CRC_OUT_2_2,II31731);
  nand NAND2_6231(WX10311,II31732,II31733);
  nand NAND2_6232(II31738,WX9692,CRC_OUT_2_1);
  nand NAND2_6233(II31739,WX9692,II31738);
  nand NAND2_6234(II31740,CRC_OUT_2_1,II31738);
  nand NAND2_6235(WX10312,II31739,II31740);
  nand NAND2_6236(II31745,WX9693,CRC_OUT_2_0);
  nand NAND2_6237(II31746,WX9693,II31745);
  nand NAND2_6238(II31747,CRC_OUT_2_0,II31745);
  nand NAND2_6239(WX10313,II31746,II31747);
  nand NAND2_6240(II34028,WX11345,WX10989);
  nand NAND2_6241(II34029,WX11345,II34028);
  nand NAND2_6242(II34030,WX10989,II34028);
  nand NAND2_6243(II34027,II34029,II34030);
  nand NAND2_6244(II34035,WX11053,II34027);
  nand NAND2_6245(II34036,WX11053,II34035);
  nand NAND2_6246(II34037,II34027,II34035);
  nand NAND2_6247(II34026,II34036,II34037);
  nand NAND2_6248(II34043,WX11117,WX11181);
  nand NAND2_6249(II34044,WX11117,II34043);
  nand NAND2_6250(II34045,WX11181,II34043);
  nand NAND2_6251(II34042,II34044,II34045);
  nand NAND2_6252(II34050,II34026,II34042);
  nand NAND2_6253(II34051,II34026,II34050);
  nand NAND2_6254(II34052,II34042,II34050);
  nand NAND2_6255(WX11244,II34051,II34052);
  nand NAND2_6256(II34059,WX11345,WX10991);
  nand NAND2_6257(II34060,WX11345,II34059);
  nand NAND2_6258(II34061,WX10991,II34059);
  nand NAND2_6259(II34058,II34060,II34061);
  nand NAND2_6260(II34066,WX11055,II34058);
  nand NAND2_6261(II34067,WX11055,II34066);
  nand NAND2_6262(II34068,II34058,II34066);
  nand NAND2_6263(II34057,II34067,II34068);
  nand NAND2_6264(II34074,WX11119,WX11183);
  nand NAND2_6265(II34075,WX11119,II34074);
  nand NAND2_6266(II34076,WX11183,II34074);
  nand NAND2_6267(II34073,II34075,II34076);
  nand NAND2_6268(II34081,II34057,II34073);
  nand NAND2_6269(II34082,II34057,II34081);
  nand NAND2_6270(II34083,II34073,II34081);
  nand NAND2_6271(WX11245,II34082,II34083);
  nand NAND2_6272(II34090,WX11345,WX10993);
  nand NAND2_6273(II34091,WX11345,II34090);
  nand NAND2_6274(II34092,WX10993,II34090);
  nand NAND2_6275(II34089,II34091,II34092);
  nand NAND2_6276(II34097,WX11057,II34089);
  nand NAND2_6277(II34098,WX11057,II34097);
  nand NAND2_6278(II34099,II34089,II34097);
  nand NAND2_6279(II34088,II34098,II34099);
  nand NAND2_6280(II34105,WX11121,WX11185);
  nand NAND2_6281(II34106,WX11121,II34105);
  nand NAND2_6282(II34107,WX11185,II34105);
  nand NAND2_6283(II34104,II34106,II34107);
  nand NAND2_6284(II34112,II34088,II34104);
  nand NAND2_6285(II34113,II34088,II34112);
  nand NAND2_6286(II34114,II34104,II34112);
  nand NAND2_6287(WX11246,II34113,II34114);
  nand NAND2_6288(II34121,WX11345,WX10995);
  nand NAND2_6289(II34122,WX11345,II34121);
  nand NAND2_6290(II34123,WX10995,II34121);
  nand NAND2_6291(II34120,II34122,II34123);
  nand NAND2_6292(II34128,WX11059,II34120);
  nand NAND2_6293(II34129,WX11059,II34128);
  nand NAND2_6294(II34130,II34120,II34128);
  nand NAND2_6295(II34119,II34129,II34130);
  nand NAND2_6296(II34136,WX11123,WX11187);
  nand NAND2_6297(II34137,WX11123,II34136);
  nand NAND2_6298(II34138,WX11187,II34136);
  nand NAND2_6299(II34135,II34137,II34138);
  nand NAND2_6300(II34143,II34119,II34135);
  nand NAND2_6301(II34144,II34119,II34143);
  nand NAND2_6302(II34145,II34135,II34143);
  nand NAND2_6303(WX11247,II34144,II34145);
  nand NAND2_6304(II34152,WX11345,WX10997);
  nand NAND2_6305(II34153,WX11345,II34152);
  nand NAND2_6306(II34154,WX10997,II34152);
  nand NAND2_6307(II34151,II34153,II34154);
  nand NAND2_6308(II34159,WX11061,II34151);
  nand NAND2_6309(II34160,WX11061,II34159);
  nand NAND2_6310(II34161,II34151,II34159);
  nand NAND2_6311(II34150,II34160,II34161);
  nand NAND2_6312(II34167,WX11125,WX11189);
  nand NAND2_6313(II34168,WX11125,II34167);
  nand NAND2_6314(II34169,WX11189,II34167);
  nand NAND2_6315(II34166,II34168,II34169);
  nand NAND2_6316(II34174,II34150,II34166);
  nand NAND2_6317(II34175,II34150,II34174);
  nand NAND2_6318(II34176,II34166,II34174);
  nand NAND2_6319(WX11248,II34175,II34176);
  nand NAND2_6320(II34183,WX11345,WX10999);
  nand NAND2_6321(II34184,WX11345,II34183);
  nand NAND2_6322(II34185,WX10999,II34183);
  nand NAND2_6323(II34182,II34184,II34185);
  nand NAND2_6324(II34190,WX11063,II34182);
  nand NAND2_6325(II34191,WX11063,II34190);
  nand NAND2_6326(II34192,II34182,II34190);
  nand NAND2_6327(II34181,II34191,II34192);
  nand NAND2_6328(II34198,WX11127,WX11191);
  nand NAND2_6329(II34199,WX11127,II34198);
  nand NAND2_6330(II34200,WX11191,II34198);
  nand NAND2_6331(II34197,II34199,II34200);
  nand NAND2_6332(II34205,II34181,II34197);
  nand NAND2_6333(II34206,II34181,II34205);
  nand NAND2_6334(II34207,II34197,II34205);
  nand NAND2_6335(WX11249,II34206,II34207);
  nand NAND2_6336(II34214,WX11345,WX11001);
  nand NAND2_6337(II34215,WX11345,II34214);
  nand NAND2_6338(II34216,WX11001,II34214);
  nand NAND2_6339(II34213,II34215,II34216);
  nand NAND2_6340(II34221,WX11065,II34213);
  nand NAND2_6341(II34222,WX11065,II34221);
  nand NAND2_6342(II34223,II34213,II34221);
  nand NAND2_6343(II34212,II34222,II34223);
  nand NAND2_6344(II34229,WX11129,WX11193);
  nand NAND2_6345(II34230,WX11129,II34229);
  nand NAND2_6346(II34231,WX11193,II34229);
  nand NAND2_6347(II34228,II34230,II34231);
  nand NAND2_6348(II34236,II34212,II34228);
  nand NAND2_6349(II34237,II34212,II34236);
  nand NAND2_6350(II34238,II34228,II34236);
  nand NAND2_6351(WX11250,II34237,II34238);
  nand NAND2_6352(II34245,WX11345,WX11003);
  nand NAND2_6353(II34246,WX11345,II34245);
  nand NAND2_6354(II34247,WX11003,II34245);
  nand NAND2_6355(II34244,II34246,II34247);
  nand NAND2_6356(II34252,WX11067,II34244);
  nand NAND2_6357(II34253,WX11067,II34252);
  nand NAND2_6358(II34254,II34244,II34252);
  nand NAND2_6359(II34243,II34253,II34254);
  nand NAND2_6360(II34260,WX11131,WX11195);
  nand NAND2_6361(II34261,WX11131,II34260);
  nand NAND2_6362(II34262,WX11195,II34260);
  nand NAND2_6363(II34259,II34261,II34262);
  nand NAND2_6364(II34267,II34243,II34259);
  nand NAND2_6365(II34268,II34243,II34267);
  nand NAND2_6366(II34269,II34259,II34267);
  nand NAND2_6367(WX11251,II34268,II34269);
  nand NAND2_6368(II34276,WX11345,WX11005);
  nand NAND2_6369(II34277,WX11345,II34276);
  nand NAND2_6370(II34278,WX11005,II34276);
  nand NAND2_6371(II34275,II34277,II34278);
  nand NAND2_6372(II34283,WX11069,II34275);
  nand NAND2_6373(II34284,WX11069,II34283);
  nand NAND2_6374(II34285,II34275,II34283);
  nand NAND2_6375(II34274,II34284,II34285);
  nand NAND2_6376(II34291,WX11133,WX11197);
  nand NAND2_6377(II34292,WX11133,II34291);
  nand NAND2_6378(II34293,WX11197,II34291);
  nand NAND2_6379(II34290,II34292,II34293);
  nand NAND2_6380(II34298,II34274,II34290);
  nand NAND2_6381(II34299,II34274,II34298);
  nand NAND2_6382(II34300,II34290,II34298);
  nand NAND2_6383(WX11252,II34299,II34300);
  nand NAND2_6384(II34307,WX11345,WX11007);
  nand NAND2_6385(II34308,WX11345,II34307);
  nand NAND2_6386(II34309,WX11007,II34307);
  nand NAND2_6387(II34306,II34308,II34309);
  nand NAND2_6388(II34314,WX11071,II34306);
  nand NAND2_6389(II34315,WX11071,II34314);
  nand NAND2_6390(II34316,II34306,II34314);
  nand NAND2_6391(II34305,II34315,II34316);
  nand NAND2_6392(II34322,WX11135,WX11199);
  nand NAND2_6393(II34323,WX11135,II34322);
  nand NAND2_6394(II34324,WX11199,II34322);
  nand NAND2_6395(II34321,II34323,II34324);
  nand NAND2_6396(II34329,II34305,II34321);
  nand NAND2_6397(II34330,II34305,II34329);
  nand NAND2_6398(II34331,II34321,II34329);
  nand NAND2_6399(WX11253,II34330,II34331);
  nand NAND2_6400(II34338,WX11345,WX11009);
  nand NAND2_6401(II34339,WX11345,II34338);
  nand NAND2_6402(II34340,WX11009,II34338);
  nand NAND2_6403(II34337,II34339,II34340);
  nand NAND2_6404(II34345,WX11073,II34337);
  nand NAND2_6405(II34346,WX11073,II34345);
  nand NAND2_6406(II34347,II34337,II34345);
  nand NAND2_6407(II34336,II34346,II34347);
  nand NAND2_6408(II34353,WX11137,WX11201);
  nand NAND2_6409(II34354,WX11137,II34353);
  nand NAND2_6410(II34355,WX11201,II34353);
  nand NAND2_6411(II34352,II34354,II34355);
  nand NAND2_6412(II34360,II34336,II34352);
  nand NAND2_6413(II34361,II34336,II34360);
  nand NAND2_6414(II34362,II34352,II34360);
  nand NAND2_6415(WX11254,II34361,II34362);
  nand NAND2_6416(II34369,WX11345,WX11011);
  nand NAND2_6417(II34370,WX11345,II34369);
  nand NAND2_6418(II34371,WX11011,II34369);
  nand NAND2_6419(II34368,II34370,II34371);
  nand NAND2_6420(II34376,WX11075,II34368);
  nand NAND2_6421(II34377,WX11075,II34376);
  nand NAND2_6422(II34378,II34368,II34376);
  nand NAND2_6423(II34367,II34377,II34378);
  nand NAND2_6424(II34384,WX11139,WX11203);
  nand NAND2_6425(II34385,WX11139,II34384);
  nand NAND2_6426(II34386,WX11203,II34384);
  nand NAND2_6427(II34383,II34385,II34386);
  nand NAND2_6428(II34391,II34367,II34383);
  nand NAND2_6429(II34392,II34367,II34391);
  nand NAND2_6430(II34393,II34383,II34391);
  nand NAND2_6431(WX11255,II34392,II34393);
  nand NAND2_6432(II34400,WX11345,WX11013);
  nand NAND2_6433(II34401,WX11345,II34400);
  nand NAND2_6434(II34402,WX11013,II34400);
  nand NAND2_6435(II34399,II34401,II34402);
  nand NAND2_6436(II34407,WX11077,II34399);
  nand NAND2_6437(II34408,WX11077,II34407);
  nand NAND2_6438(II34409,II34399,II34407);
  nand NAND2_6439(II34398,II34408,II34409);
  nand NAND2_6440(II34415,WX11141,WX11205);
  nand NAND2_6441(II34416,WX11141,II34415);
  nand NAND2_6442(II34417,WX11205,II34415);
  nand NAND2_6443(II34414,II34416,II34417);
  nand NAND2_6444(II34422,II34398,II34414);
  nand NAND2_6445(II34423,II34398,II34422);
  nand NAND2_6446(II34424,II34414,II34422);
  nand NAND2_6447(WX11256,II34423,II34424);
  nand NAND2_6448(II34431,WX11345,WX11015);
  nand NAND2_6449(II34432,WX11345,II34431);
  nand NAND2_6450(II34433,WX11015,II34431);
  nand NAND2_6451(II34430,II34432,II34433);
  nand NAND2_6452(II34438,WX11079,II34430);
  nand NAND2_6453(II34439,WX11079,II34438);
  nand NAND2_6454(II34440,II34430,II34438);
  nand NAND2_6455(II34429,II34439,II34440);
  nand NAND2_6456(II34446,WX11143,WX11207);
  nand NAND2_6457(II34447,WX11143,II34446);
  nand NAND2_6458(II34448,WX11207,II34446);
  nand NAND2_6459(II34445,II34447,II34448);
  nand NAND2_6460(II34453,II34429,II34445);
  nand NAND2_6461(II34454,II34429,II34453);
  nand NAND2_6462(II34455,II34445,II34453);
  nand NAND2_6463(WX11257,II34454,II34455);
  nand NAND2_6464(II34462,WX11345,WX11017);
  nand NAND2_6465(II34463,WX11345,II34462);
  nand NAND2_6466(II34464,WX11017,II34462);
  nand NAND2_6467(II34461,II34463,II34464);
  nand NAND2_6468(II34469,WX11081,II34461);
  nand NAND2_6469(II34470,WX11081,II34469);
  nand NAND2_6470(II34471,II34461,II34469);
  nand NAND2_6471(II34460,II34470,II34471);
  nand NAND2_6472(II34477,WX11145,WX11209);
  nand NAND2_6473(II34478,WX11145,II34477);
  nand NAND2_6474(II34479,WX11209,II34477);
  nand NAND2_6475(II34476,II34478,II34479);
  nand NAND2_6476(II34484,II34460,II34476);
  nand NAND2_6477(II34485,II34460,II34484);
  nand NAND2_6478(II34486,II34476,II34484);
  nand NAND2_6479(WX11258,II34485,II34486);
  nand NAND2_6480(II34493,WX11345,WX11019);
  nand NAND2_6481(II34494,WX11345,II34493);
  nand NAND2_6482(II34495,WX11019,II34493);
  nand NAND2_6483(II34492,II34494,II34495);
  nand NAND2_6484(II34500,WX11083,II34492);
  nand NAND2_6485(II34501,WX11083,II34500);
  nand NAND2_6486(II34502,II34492,II34500);
  nand NAND2_6487(II34491,II34501,II34502);
  nand NAND2_6488(II34508,WX11147,WX11211);
  nand NAND2_6489(II34509,WX11147,II34508);
  nand NAND2_6490(II34510,WX11211,II34508);
  nand NAND2_6491(II34507,II34509,II34510);
  nand NAND2_6492(II34515,II34491,II34507);
  nand NAND2_6493(II34516,II34491,II34515);
  nand NAND2_6494(II34517,II34507,II34515);
  nand NAND2_6495(WX11259,II34516,II34517);
  nand NAND2_6496(II34524,WX11346,WX11021);
  nand NAND2_6497(II34525,WX11346,II34524);
  nand NAND2_6498(II34526,WX11021,II34524);
  nand NAND2_6499(II34523,II34525,II34526);
  nand NAND2_6500(II34531,WX11085,II34523);
  nand NAND2_6501(II34532,WX11085,II34531);
  nand NAND2_6502(II34533,II34523,II34531);
  nand NAND2_6503(II34522,II34532,II34533);
  nand NAND2_6504(II34539,WX11149,WX11213);
  nand NAND2_6505(II34540,WX11149,II34539);
  nand NAND2_6506(II34541,WX11213,II34539);
  nand NAND2_6507(II34538,II34540,II34541);
  nand NAND2_6508(II34546,II34522,II34538);
  nand NAND2_6509(II34547,II34522,II34546);
  nand NAND2_6510(II34548,II34538,II34546);
  nand NAND2_6511(WX11260,II34547,II34548);
  nand NAND2_6512(II34555,WX11346,WX11023);
  nand NAND2_6513(II34556,WX11346,II34555);
  nand NAND2_6514(II34557,WX11023,II34555);
  nand NAND2_6515(II34554,II34556,II34557);
  nand NAND2_6516(II34562,WX11087,II34554);
  nand NAND2_6517(II34563,WX11087,II34562);
  nand NAND2_6518(II34564,II34554,II34562);
  nand NAND2_6519(II34553,II34563,II34564);
  nand NAND2_6520(II34570,WX11151,WX11215);
  nand NAND2_6521(II34571,WX11151,II34570);
  nand NAND2_6522(II34572,WX11215,II34570);
  nand NAND2_6523(II34569,II34571,II34572);
  nand NAND2_6524(II34577,II34553,II34569);
  nand NAND2_6525(II34578,II34553,II34577);
  nand NAND2_6526(II34579,II34569,II34577);
  nand NAND2_6527(WX11261,II34578,II34579);
  nand NAND2_6528(II34586,WX11346,WX11025);
  nand NAND2_6529(II34587,WX11346,II34586);
  nand NAND2_6530(II34588,WX11025,II34586);
  nand NAND2_6531(II34585,II34587,II34588);
  nand NAND2_6532(II34593,WX11089,II34585);
  nand NAND2_6533(II34594,WX11089,II34593);
  nand NAND2_6534(II34595,II34585,II34593);
  nand NAND2_6535(II34584,II34594,II34595);
  nand NAND2_6536(II34601,WX11153,WX11217);
  nand NAND2_6537(II34602,WX11153,II34601);
  nand NAND2_6538(II34603,WX11217,II34601);
  nand NAND2_6539(II34600,II34602,II34603);
  nand NAND2_6540(II34608,II34584,II34600);
  nand NAND2_6541(II34609,II34584,II34608);
  nand NAND2_6542(II34610,II34600,II34608);
  nand NAND2_6543(WX11262,II34609,II34610);
  nand NAND2_6544(II34617,WX11346,WX11027);
  nand NAND2_6545(II34618,WX11346,II34617);
  nand NAND2_6546(II34619,WX11027,II34617);
  nand NAND2_6547(II34616,II34618,II34619);
  nand NAND2_6548(II34624,WX11091,II34616);
  nand NAND2_6549(II34625,WX11091,II34624);
  nand NAND2_6550(II34626,II34616,II34624);
  nand NAND2_6551(II34615,II34625,II34626);
  nand NAND2_6552(II34632,WX11155,WX11219);
  nand NAND2_6553(II34633,WX11155,II34632);
  nand NAND2_6554(II34634,WX11219,II34632);
  nand NAND2_6555(II34631,II34633,II34634);
  nand NAND2_6556(II34639,II34615,II34631);
  nand NAND2_6557(II34640,II34615,II34639);
  nand NAND2_6558(II34641,II34631,II34639);
  nand NAND2_6559(WX11263,II34640,II34641);
  nand NAND2_6560(II34648,WX11346,WX11029);
  nand NAND2_6561(II34649,WX11346,II34648);
  nand NAND2_6562(II34650,WX11029,II34648);
  nand NAND2_6563(II34647,II34649,II34650);
  nand NAND2_6564(II34655,WX11093,II34647);
  nand NAND2_6565(II34656,WX11093,II34655);
  nand NAND2_6566(II34657,II34647,II34655);
  nand NAND2_6567(II34646,II34656,II34657);
  nand NAND2_6568(II34663,WX11157,WX11221);
  nand NAND2_6569(II34664,WX11157,II34663);
  nand NAND2_6570(II34665,WX11221,II34663);
  nand NAND2_6571(II34662,II34664,II34665);
  nand NAND2_6572(II34670,II34646,II34662);
  nand NAND2_6573(II34671,II34646,II34670);
  nand NAND2_6574(II34672,II34662,II34670);
  nand NAND2_6575(WX11264,II34671,II34672);
  nand NAND2_6576(II34679,WX11346,WX11031);
  nand NAND2_6577(II34680,WX11346,II34679);
  nand NAND2_6578(II34681,WX11031,II34679);
  nand NAND2_6579(II34678,II34680,II34681);
  nand NAND2_6580(II34686,WX11095,II34678);
  nand NAND2_6581(II34687,WX11095,II34686);
  nand NAND2_6582(II34688,II34678,II34686);
  nand NAND2_6583(II34677,II34687,II34688);
  nand NAND2_6584(II34694,WX11159,WX11223);
  nand NAND2_6585(II34695,WX11159,II34694);
  nand NAND2_6586(II34696,WX11223,II34694);
  nand NAND2_6587(II34693,II34695,II34696);
  nand NAND2_6588(II34701,II34677,II34693);
  nand NAND2_6589(II34702,II34677,II34701);
  nand NAND2_6590(II34703,II34693,II34701);
  nand NAND2_6591(WX11265,II34702,II34703);
  nand NAND2_6592(II34710,WX11346,WX11033);
  nand NAND2_6593(II34711,WX11346,II34710);
  nand NAND2_6594(II34712,WX11033,II34710);
  nand NAND2_6595(II34709,II34711,II34712);
  nand NAND2_6596(II34717,WX11097,II34709);
  nand NAND2_6597(II34718,WX11097,II34717);
  nand NAND2_6598(II34719,II34709,II34717);
  nand NAND2_6599(II34708,II34718,II34719);
  nand NAND2_6600(II34725,WX11161,WX11225);
  nand NAND2_6601(II34726,WX11161,II34725);
  nand NAND2_6602(II34727,WX11225,II34725);
  nand NAND2_6603(II34724,II34726,II34727);
  nand NAND2_6604(II34732,II34708,II34724);
  nand NAND2_6605(II34733,II34708,II34732);
  nand NAND2_6606(II34734,II34724,II34732);
  nand NAND2_6607(WX11266,II34733,II34734);
  nand NAND2_6608(II34741,WX11346,WX11035);
  nand NAND2_6609(II34742,WX11346,II34741);
  nand NAND2_6610(II34743,WX11035,II34741);
  nand NAND2_6611(II34740,II34742,II34743);
  nand NAND2_6612(II34748,WX11099,II34740);
  nand NAND2_6613(II34749,WX11099,II34748);
  nand NAND2_6614(II34750,II34740,II34748);
  nand NAND2_6615(II34739,II34749,II34750);
  nand NAND2_6616(II34756,WX11163,WX11227);
  nand NAND2_6617(II34757,WX11163,II34756);
  nand NAND2_6618(II34758,WX11227,II34756);
  nand NAND2_6619(II34755,II34757,II34758);
  nand NAND2_6620(II34763,II34739,II34755);
  nand NAND2_6621(II34764,II34739,II34763);
  nand NAND2_6622(II34765,II34755,II34763);
  nand NAND2_6623(WX11267,II34764,II34765);
  nand NAND2_6624(II34772,WX11346,WX11037);
  nand NAND2_6625(II34773,WX11346,II34772);
  nand NAND2_6626(II34774,WX11037,II34772);
  nand NAND2_6627(II34771,II34773,II34774);
  nand NAND2_6628(II34779,WX11101,II34771);
  nand NAND2_6629(II34780,WX11101,II34779);
  nand NAND2_6630(II34781,II34771,II34779);
  nand NAND2_6631(II34770,II34780,II34781);
  nand NAND2_6632(II34787,WX11165,WX11229);
  nand NAND2_6633(II34788,WX11165,II34787);
  nand NAND2_6634(II34789,WX11229,II34787);
  nand NAND2_6635(II34786,II34788,II34789);
  nand NAND2_6636(II34794,II34770,II34786);
  nand NAND2_6637(II34795,II34770,II34794);
  nand NAND2_6638(II34796,II34786,II34794);
  nand NAND2_6639(WX11268,II34795,II34796);
  nand NAND2_6640(II34803,WX11346,WX11039);
  nand NAND2_6641(II34804,WX11346,II34803);
  nand NAND2_6642(II34805,WX11039,II34803);
  nand NAND2_6643(II34802,II34804,II34805);
  nand NAND2_6644(II34810,WX11103,II34802);
  nand NAND2_6645(II34811,WX11103,II34810);
  nand NAND2_6646(II34812,II34802,II34810);
  nand NAND2_6647(II34801,II34811,II34812);
  nand NAND2_6648(II34818,WX11167,WX11231);
  nand NAND2_6649(II34819,WX11167,II34818);
  nand NAND2_6650(II34820,WX11231,II34818);
  nand NAND2_6651(II34817,II34819,II34820);
  nand NAND2_6652(II34825,II34801,II34817);
  nand NAND2_6653(II34826,II34801,II34825);
  nand NAND2_6654(II34827,II34817,II34825);
  nand NAND2_6655(WX11269,II34826,II34827);
  nand NAND2_6656(II34834,WX11346,WX11041);
  nand NAND2_6657(II34835,WX11346,II34834);
  nand NAND2_6658(II34836,WX11041,II34834);
  nand NAND2_6659(II34833,II34835,II34836);
  nand NAND2_6660(II34841,WX11105,II34833);
  nand NAND2_6661(II34842,WX11105,II34841);
  nand NAND2_6662(II34843,II34833,II34841);
  nand NAND2_6663(II34832,II34842,II34843);
  nand NAND2_6664(II34849,WX11169,WX11233);
  nand NAND2_6665(II34850,WX11169,II34849);
  nand NAND2_6666(II34851,WX11233,II34849);
  nand NAND2_6667(II34848,II34850,II34851);
  nand NAND2_6668(II34856,II34832,II34848);
  nand NAND2_6669(II34857,II34832,II34856);
  nand NAND2_6670(II34858,II34848,II34856);
  nand NAND2_6671(WX11270,II34857,II34858);
  nand NAND2_6672(II34865,WX11346,WX11043);
  nand NAND2_6673(II34866,WX11346,II34865);
  nand NAND2_6674(II34867,WX11043,II34865);
  nand NAND2_6675(II34864,II34866,II34867);
  nand NAND2_6676(II34872,WX11107,II34864);
  nand NAND2_6677(II34873,WX11107,II34872);
  nand NAND2_6678(II34874,II34864,II34872);
  nand NAND2_6679(II34863,II34873,II34874);
  nand NAND2_6680(II34880,WX11171,WX11235);
  nand NAND2_6681(II34881,WX11171,II34880);
  nand NAND2_6682(II34882,WX11235,II34880);
  nand NAND2_6683(II34879,II34881,II34882);
  nand NAND2_6684(II34887,II34863,II34879);
  nand NAND2_6685(II34888,II34863,II34887);
  nand NAND2_6686(II34889,II34879,II34887);
  nand NAND2_6687(WX11271,II34888,II34889);
  nand NAND2_6688(II34896,WX11346,WX11045);
  nand NAND2_6689(II34897,WX11346,II34896);
  nand NAND2_6690(II34898,WX11045,II34896);
  nand NAND2_6691(II34895,II34897,II34898);
  nand NAND2_6692(II34903,WX11109,II34895);
  nand NAND2_6693(II34904,WX11109,II34903);
  nand NAND2_6694(II34905,II34895,II34903);
  nand NAND2_6695(II34894,II34904,II34905);
  nand NAND2_6696(II34911,WX11173,WX11237);
  nand NAND2_6697(II34912,WX11173,II34911);
  nand NAND2_6698(II34913,WX11237,II34911);
  nand NAND2_6699(II34910,II34912,II34913);
  nand NAND2_6700(II34918,II34894,II34910);
  nand NAND2_6701(II34919,II34894,II34918);
  nand NAND2_6702(II34920,II34910,II34918);
  nand NAND2_6703(WX11272,II34919,II34920);
  nand NAND2_6704(II34927,WX11346,WX11047);
  nand NAND2_6705(II34928,WX11346,II34927);
  nand NAND2_6706(II34929,WX11047,II34927);
  nand NAND2_6707(II34926,II34928,II34929);
  nand NAND2_6708(II34934,WX11111,II34926);
  nand NAND2_6709(II34935,WX11111,II34934);
  nand NAND2_6710(II34936,II34926,II34934);
  nand NAND2_6711(II34925,II34935,II34936);
  nand NAND2_6712(II34942,WX11175,WX11239);
  nand NAND2_6713(II34943,WX11175,II34942);
  nand NAND2_6714(II34944,WX11239,II34942);
  nand NAND2_6715(II34941,II34943,II34944);
  nand NAND2_6716(II34949,II34925,II34941);
  nand NAND2_6717(II34950,II34925,II34949);
  nand NAND2_6718(II34951,II34941,II34949);
  nand NAND2_6719(WX11273,II34950,II34951);
  nand NAND2_6720(II34958,WX11346,WX11049);
  nand NAND2_6721(II34959,WX11346,II34958);
  nand NAND2_6722(II34960,WX11049,II34958);
  nand NAND2_6723(II34957,II34959,II34960);
  nand NAND2_6724(II34965,WX11113,II34957);
  nand NAND2_6725(II34966,WX11113,II34965);
  nand NAND2_6726(II34967,II34957,II34965);
  nand NAND2_6727(II34956,II34966,II34967);
  nand NAND2_6728(II34973,WX11177,WX11241);
  nand NAND2_6729(II34974,WX11177,II34973);
  nand NAND2_6730(II34975,WX11241,II34973);
  nand NAND2_6731(II34972,II34974,II34975);
  nand NAND2_6732(II34980,II34956,II34972);
  nand NAND2_6733(II34981,II34956,II34980);
  nand NAND2_6734(II34982,II34972,II34980);
  nand NAND2_6735(WX11274,II34981,II34982);
  nand NAND2_6736(II34989,WX11346,WX11051);
  nand NAND2_6737(II34990,WX11346,II34989);
  nand NAND2_6738(II34991,WX11051,II34989);
  nand NAND2_6739(II34988,II34990,II34991);
  nand NAND2_6740(II34996,WX11115,II34988);
  nand NAND2_6741(II34997,WX11115,II34996);
  nand NAND2_6742(II34998,II34988,II34996);
  nand NAND2_6743(II34987,II34997,II34998);
  nand NAND2_6744(II35004,WX11179,WX11243);
  nand NAND2_6745(II35005,WX11179,II35004);
  nand NAND2_6746(II35006,WX11243,II35004);
  nand NAND2_6747(II35003,II35005,II35006);
  nand NAND2_6748(II35011,II34987,II35003);
  nand NAND2_6749(II35012,II34987,II35011);
  nand NAND2_6750(II35013,II35003,II35011);
  nand NAND2_6751(WX11275,II35012,II35013);
  nand NAND2_6752(II35092,WX10924,WX10829);
  nand NAND2_6753(II35093,WX10924,II35092);
  nand NAND2_6754(II35094,WX10829,II35092);
  nand NAND2_6755(WX11350,II35093,II35094);
  nand NAND2_6756(II35105,WX10925,WX10831);
  nand NAND2_6757(II35106,WX10925,II35105);
  nand NAND2_6758(II35107,WX10831,II35105);
  nand NAND2_6759(WX11357,II35106,II35107);
  nand NAND2_6760(II35118,WX10926,WX10833);
  nand NAND2_6761(II35119,WX10926,II35118);
  nand NAND2_6762(II35120,WX10833,II35118);
  nand NAND2_6763(WX11364,II35119,II35120);
  nand NAND2_6764(II35131,WX10927,WX10835);
  nand NAND2_6765(II35132,WX10927,II35131);
  nand NAND2_6766(II35133,WX10835,II35131);
  nand NAND2_6767(WX11371,II35132,II35133);
  nand NAND2_6768(II35144,WX10928,WX10837);
  nand NAND2_6769(II35145,WX10928,II35144);
  nand NAND2_6770(II35146,WX10837,II35144);
  nand NAND2_6771(WX11378,II35145,II35146);
  nand NAND2_6772(II35157,WX10929,WX10839);
  nand NAND2_6773(II35158,WX10929,II35157);
  nand NAND2_6774(II35159,WX10839,II35157);
  nand NAND2_6775(WX11385,II35158,II35159);
  nand NAND2_6776(II35170,WX10930,WX10841);
  nand NAND2_6777(II35171,WX10930,II35170);
  nand NAND2_6778(II35172,WX10841,II35170);
  nand NAND2_6779(WX11392,II35171,II35172);
  nand NAND2_6780(II35183,WX10931,WX10843);
  nand NAND2_6781(II35184,WX10931,II35183);
  nand NAND2_6782(II35185,WX10843,II35183);
  nand NAND2_6783(WX11399,II35184,II35185);
  nand NAND2_6784(II35196,WX10932,WX10845);
  nand NAND2_6785(II35197,WX10932,II35196);
  nand NAND2_6786(II35198,WX10845,II35196);
  nand NAND2_6787(WX11406,II35197,II35198);
  nand NAND2_6788(II35209,WX10933,WX10847);
  nand NAND2_6789(II35210,WX10933,II35209);
  nand NAND2_6790(II35211,WX10847,II35209);
  nand NAND2_6791(WX11413,II35210,II35211);
  nand NAND2_6792(II35222,WX10934,WX10849);
  nand NAND2_6793(II35223,WX10934,II35222);
  nand NAND2_6794(II35224,WX10849,II35222);
  nand NAND2_6795(WX11420,II35223,II35224);
  nand NAND2_6796(II35235,WX10935,WX10851);
  nand NAND2_6797(II35236,WX10935,II35235);
  nand NAND2_6798(II35237,WX10851,II35235);
  nand NAND2_6799(WX11427,II35236,II35237);
  nand NAND2_6800(II35248,WX10936,WX10853);
  nand NAND2_6801(II35249,WX10936,II35248);
  nand NAND2_6802(II35250,WX10853,II35248);
  nand NAND2_6803(WX11434,II35249,II35250);
  nand NAND2_6804(II35261,WX10937,WX10855);
  nand NAND2_6805(II35262,WX10937,II35261);
  nand NAND2_6806(II35263,WX10855,II35261);
  nand NAND2_6807(WX11441,II35262,II35263);
  nand NAND2_6808(II35274,WX10938,WX10857);
  nand NAND2_6809(II35275,WX10938,II35274);
  nand NAND2_6810(II35276,WX10857,II35274);
  nand NAND2_6811(WX11448,II35275,II35276);
  nand NAND2_6812(II35287,WX10939,WX10859);
  nand NAND2_6813(II35288,WX10939,II35287);
  nand NAND2_6814(II35289,WX10859,II35287);
  nand NAND2_6815(WX11455,II35288,II35289);
  nand NAND2_6816(II35300,WX10940,WX10861);
  nand NAND2_6817(II35301,WX10940,II35300);
  nand NAND2_6818(II35302,WX10861,II35300);
  nand NAND2_6819(WX11462,II35301,II35302);
  nand NAND2_6820(II35313,WX10941,WX10863);
  nand NAND2_6821(II35314,WX10941,II35313);
  nand NAND2_6822(II35315,WX10863,II35313);
  nand NAND2_6823(WX11469,II35314,II35315);
  nand NAND2_6824(II35326,WX10942,WX10865);
  nand NAND2_6825(II35327,WX10942,II35326);
  nand NAND2_6826(II35328,WX10865,II35326);
  nand NAND2_6827(WX11476,II35327,II35328);
  nand NAND2_6828(II35339,WX10943,WX10867);
  nand NAND2_6829(II35340,WX10943,II35339);
  nand NAND2_6830(II35341,WX10867,II35339);
  nand NAND2_6831(WX11483,II35340,II35341);
  nand NAND2_6832(II35352,WX10944,WX10869);
  nand NAND2_6833(II35353,WX10944,II35352);
  nand NAND2_6834(II35354,WX10869,II35352);
  nand NAND2_6835(WX11490,II35353,II35354);
  nand NAND2_6836(II35365,WX10945,WX10871);
  nand NAND2_6837(II35366,WX10945,II35365);
  nand NAND2_6838(II35367,WX10871,II35365);
  nand NAND2_6839(WX11497,II35366,II35367);
  nand NAND2_6840(II35378,WX10946,WX10873);
  nand NAND2_6841(II35379,WX10946,II35378);
  nand NAND2_6842(II35380,WX10873,II35378);
  nand NAND2_6843(WX11504,II35379,II35380);
  nand NAND2_6844(II35391,WX10947,WX10875);
  nand NAND2_6845(II35392,WX10947,II35391);
  nand NAND2_6846(II35393,WX10875,II35391);
  nand NAND2_6847(WX11511,II35392,II35393);
  nand NAND2_6848(II35404,WX10948,WX10877);
  nand NAND2_6849(II35405,WX10948,II35404);
  nand NAND2_6850(II35406,WX10877,II35404);
  nand NAND2_6851(WX11518,II35405,II35406);
  nand NAND2_6852(II35417,WX10949,WX10879);
  nand NAND2_6853(II35418,WX10949,II35417);
  nand NAND2_6854(II35419,WX10879,II35417);
  nand NAND2_6855(WX11525,II35418,II35419);
  nand NAND2_6856(II35430,WX10950,WX10881);
  nand NAND2_6857(II35431,WX10950,II35430);
  nand NAND2_6858(II35432,WX10881,II35430);
  nand NAND2_6859(WX11532,II35431,II35432);
  nand NAND2_6860(II35443,WX10951,WX10883);
  nand NAND2_6861(II35444,WX10951,II35443);
  nand NAND2_6862(II35445,WX10883,II35443);
  nand NAND2_6863(WX11539,II35444,II35445);
  nand NAND2_6864(II35456,WX10952,WX10885);
  nand NAND2_6865(II35457,WX10952,II35456);
  nand NAND2_6866(II35458,WX10885,II35456);
  nand NAND2_6867(WX11546,II35457,II35458);
  nand NAND2_6868(II35469,WX10953,WX10887);
  nand NAND2_6869(II35470,WX10953,II35469);
  nand NAND2_6870(II35471,WX10887,II35469);
  nand NAND2_6871(WX11553,II35470,II35471);
  nand NAND2_6872(II35482,WX10954,WX10889);
  nand NAND2_6873(II35483,WX10954,II35482);
  nand NAND2_6874(II35484,WX10889,II35482);
  nand NAND2_6875(WX11560,II35483,II35484);
  nand NAND2_6876(II35495,WX10955,WX10891);
  nand NAND2_6877(II35496,WX10955,II35495);
  nand NAND2_6878(II35497,WX10891,II35495);
  nand NAND2_6879(WX11567,II35496,II35497);
  nand NAND2_6880(II35510,WX10971,CRC_OUT_1_31);
  nand NAND2_6881(II35511,WX10971,II35510);
  nand NAND2_6882(II35512,CRC_OUT_1_31,II35510);
  nand NAND2_6883(II35509,II35511,II35512);
  nand NAND2_6884(II35517,CRC_OUT_1_15,II35509);
  nand NAND2_6885(II35518,CRC_OUT_1_15,II35517);
  nand NAND2_6886(II35519,II35509,II35517);
  nand NAND2_6887(WX11575,II35518,II35519);
  nand NAND2_6888(II35525,WX10976,CRC_OUT_1_31);
  nand NAND2_6889(II35526,WX10976,II35525);
  nand NAND2_6890(II35527,CRC_OUT_1_31,II35525);
  nand NAND2_6891(II35524,II35526,II35527);
  nand NAND2_6892(II35532,CRC_OUT_1_10,II35524);
  nand NAND2_6893(II35533,CRC_OUT_1_10,II35532);
  nand NAND2_6894(II35534,II35524,II35532);
  nand NAND2_6895(WX11576,II35533,II35534);
  nand NAND2_6896(II35540,WX10983,CRC_OUT_1_31);
  nand NAND2_6897(II35541,WX10983,II35540);
  nand NAND2_6898(II35542,CRC_OUT_1_31,II35540);
  nand NAND2_6899(II35539,II35541,II35542);
  nand NAND2_6900(II35547,CRC_OUT_1_3,II35539);
  nand NAND2_6901(II35548,CRC_OUT_1_3,II35547);
  nand NAND2_6902(II35549,II35539,II35547);
  nand NAND2_6903(WX11577,II35548,II35549);
  nand NAND2_6904(II35554,WX10987,CRC_OUT_1_31);
  nand NAND2_6905(II35555,WX10987,II35554);
  nand NAND2_6906(II35556,CRC_OUT_1_31,II35554);
  nand NAND2_6907(WX11578,II35555,II35556);
  nand NAND2_6908(II35561,WX10956,CRC_OUT_1_30);
  nand NAND2_6909(II35562,WX10956,II35561);
  nand NAND2_6910(II35563,CRC_OUT_1_30,II35561);
  nand NAND2_6911(WX11579,II35562,II35563);
  nand NAND2_6912(II35568,WX10957,CRC_OUT_1_29);
  nand NAND2_6913(II35569,WX10957,II35568);
  nand NAND2_6914(II35570,CRC_OUT_1_29,II35568);
  nand NAND2_6915(WX11580,II35569,II35570);
  nand NAND2_6916(II35575,WX10958,CRC_OUT_1_28);
  nand NAND2_6917(II35576,WX10958,II35575);
  nand NAND2_6918(II35577,CRC_OUT_1_28,II35575);
  nand NAND2_6919(WX11581,II35576,II35577);
  nand NAND2_6920(II35582,WX10959,CRC_OUT_1_27);
  nand NAND2_6921(II35583,WX10959,II35582);
  nand NAND2_6922(II35584,CRC_OUT_1_27,II35582);
  nand NAND2_6923(WX11582,II35583,II35584);
  nand NAND2_6924(II35589,WX10960,CRC_OUT_1_26);
  nand NAND2_6925(II35590,WX10960,II35589);
  nand NAND2_6926(II35591,CRC_OUT_1_26,II35589);
  nand NAND2_6927(WX11583,II35590,II35591);
  nand NAND2_6928(II35596,WX10961,CRC_OUT_1_25);
  nand NAND2_6929(II35597,WX10961,II35596);
  nand NAND2_6930(II35598,CRC_OUT_1_25,II35596);
  nand NAND2_6931(WX11584,II35597,II35598);
  nand NAND2_6932(II35603,WX10962,CRC_OUT_1_24);
  nand NAND2_6933(II35604,WX10962,II35603);
  nand NAND2_6934(II35605,CRC_OUT_1_24,II35603);
  nand NAND2_6935(WX11585,II35604,II35605);
  nand NAND2_6936(II35610,WX10963,CRC_OUT_1_23);
  nand NAND2_6937(II35611,WX10963,II35610);
  nand NAND2_6938(II35612,CRC_OUT_1_23,II35610);
  nand NAND2_6939(WX11586,II35611,II35612);
  nand NAND2_6940(II35617,WX10964,CRC_OUT_1_22);
  nand NAND2_6941(II35618,WX10964,II35617);
  nand NAND2_6942(II35619,CRC_OUT_1_22,II35617);
  nand NAND2_6943(WX11587,II35618,II35619);
  nand NAND2_6944(II35624,WX10965,CRC_OUT_1_21);
  nand NAND2_6945(II35625,WX10965,II35624);
  nand NAND2_6946(II35626,CRC_OUT_1_21,II35624);
  nand NAND2_6947(WX11588,II35625,II35626);
  nand NAND2_6948(II35631,WX10966,CRC_OUT_1_20);
  nand NAND2_6949(II35632,WX10966,II35631);
  nand NAND2_6950(II35633,CRC_OUT_1_20,II35631);
  nand NAND2_6951(WX11589,II35632,II35633);
  nand NAND2_6952(II35638,WX10967,CRC_OUT_1_19);
  nand NAND2_6953(II35639,WX10967,II35638);
  nand NAND2_6954(II35640,CRC_OUT_1_19,II35638);
  nand NAND2_6955(WX11590,II35639,II35640);
  nand NAND2_6956(II35645,WX10968,CRC_OUT_1_18);
  nand NAND2_6957(II35646,WX10968,II35645);
  nand NAND2_6958(II35647,CRC_OUT_1_18,II35645);
  nand NAND2_6959(WX11591,II35646,II35647);
  nand NAND2_6960(II35652,WX10969,CRC_OUT_1_17);
  nand NAND2_6961(II35653,WX10969,II35652);
  nand NAND2_6962(II35654,CRC_OUT_1_17,II35652);
  nand NAND2_6963(WX11592,II35653,II35654);
  nand NAND2_6964(II35659,WX10970,CRC_OUT_1_16);
  nand NAND2_6965(II35660,WX10970,II35659);
  nand NAND2_6966(II35661,CRC_OUT_1_16,II35659);
  nand NAND2_6967(WX11593,II35660,II35661);
  nand NAND2_6968(II35666,WX10972,CRC_OUT_1_14);
  nand NAND2_6969(II35667,WX10972,II35666);
  nand NAND2_6970(II35668,CRC_OUT_1_14,II35666);
  nand NAND2_6971(WX11594,II35667,II35668);
  nand NAND2_6972(II35673,WX10973,CRC_OUT_1_13);
  nand NAND2_6973(II35674,WX10973,II35673);
  nand NAND2_6974(II35675,CRC_OUT_1_13,II35673);
  nand NAND2_6975(WX11595,II35674,II35675);
  nand NAND2_6976(II35680,WX10974,CRC_OUT_1_12);
  nand NAND2_6977(II35681,WX10974,II35680);
  nand NAND2_6978(II35682,CRC_OUT_1_12,II35680);
  nand NAND2_6979(WX11596,II35681,II35682);
  nand NAND2_6980(II35687,WX10975,CRC_OUT_1_11);
  nand NAND2_6981(II35688,WX10975,II35687);
  nand NAND2_6982(II35689,CRC_OUT_1_11,II35687);
  nand NAND2_6983(WX11597,II35688,II35689);
  nand NAND2_6984(II35694,WX10977,CRC_OUT_1_9);
  nand NAND2_6985(II35695,WX10977,II35694);
  nand NAND2_6986(II35696,CRC_OUT_1_9,II35694);
  nand NAND2_6987(WX11598,II35695,II35696);
  nand NAND2_6988(II35701,WX10978,CRC_OUT_1_8);
  nand NAND2_6989(II35702,WX10978,II35701);
  nand NAND2_6990(II35703,CRC_OUT_1_8,II35701);
  nand NAND2_6991(WX11599,II35702,II35703);
  nand NAND2_6992(II35708,WX10979,CRC_OUT_1_7);
  nand NAND2_6993(II35709,WX10979,II35708);
  nand NAND2_6994(II35710,CRC_OUT_1_7,II35708);
  nand NAND2_6995(WX11600,II35709,II35710);
  nand NAND2_6996(II35715,WX10980,CRC_OUT_1_6);
  nand NAND2_6997(II35716,WX10980,II35715);
  nand NAND2_6998(II35717,CRC_OUT_1_6,II35715);
  nand NAND2_6999(WX11601,II35716,II35717);
  nand NAND2_7000(II35722,WX10981,CRC_OUT_1_5);
  nand NAND2_7001(II35723,WX10981,II35722);
  nand NAND2_7002(II35724,CRC_OUT_1_5,II35722);
  nand NAND2_7003(WX11602,II35723,II35724);
  nand NAND2_7004(II35729,WX10982,CRC_OUT_1_4);
  nand NAND2_7005(II35730,WX10982,II35729);
  nand NAND2_7006(II35731,CRC_OUT_1_4,II35729);
  nand NAND2_7007(WX11603,II35730,II35731);
  nand NAND2_7008(II35736,WX10984,CRC_OUT_1_2);
  nand NAND2_7009(II35737,WX10984,II35736);
  nand NAND2_7010(II35738,CRC_OUT_1_2,II35736);
  nand NAND2_7011(WX11604,II35737,II35738);
  nand NAND2_7012(II35743,WX10985,CRC_OUT_1_1);
  nand NAND2_7013(II35744,WX10985,II35743);
  nand NAND2_7014(II35745,CRC_OUT_1_1,II35743);
  nand NAND2_7015(WX11605,II35744,II35745);
  nand NAND2_7016(II35750,WX10986,CRC_OUT_1_0);
  nand NAND2_7017(II35751,WX10986,II35750);
  nand NAND2_7018(II35752,CRC_OUT_1_0,II35750);
  nand NAND2_7019(WX11606,II35751,II35752);

endmodule