module apex7(CAPSD, CAT0, CAT1, CAT2, CAT3, CAT4, CAT5, VACC, MMERR, IBT0, IBT1, IBT2, ICLR, LSD, ACCRPY, VERR_N, RATR, MARSSR, VLENESR, VSUMESR, PLUTO0, PLUTO1, PLUTO2, PLUTO3, PLUTO4, PLUTO5, ORWD_N, OWL_N, PY, \END , FBI, WATCH, OVACC, KBG_N, DEL1, COMPPAR, VST0, VST1, STAR0, STAR1, STAR2, STAR3, BULL0, BULL1, BULL2, BULL3, BULL4, BULL5, BULL6, SDO, LSD_P, ACCRPY_P, VERR_F, RATR_P, MARSSR_P, VLENESR_P, VSUMESR_P, PLUTO0_P, PLUTO1_P, PLUTO2_P, PLUTO3_P, PLUTO4_P, PLUTO5_P, ORWD_F, OWL_F, PY_P, END_P, FBI_P, WATCH_P, OVACC_P, KBG_F, DEL1_P, COMPPAR_P, VST0_P, VST1_P, STAR0_P, STAR1_P, STAR2_P, STAR3_P, BULL0_P, BULL1_P, BULL2_P, BULL3_P, BULL4_P, BULL5_P, BULL6_P);
input
  PLUTO0,
  PLUTO1,
  PLUTO2,
  PLUTO3,
  PLUTO4,
  PLUTO5,
  PY,
  VST0,
  VST1,
  VLENESR,
  BULL0,
  BULL1,
  BULL2,
  BULL3,
  BULL4,
  BULL5,
  BULL6,
  MMERR,
  VERR_N,
  MARSSR,
  \END ,
  WATCH,
  FBI,
  STAR0,
  STAR1,
  STAR2,
  STAR3,
  ACCRPY,
  IBT0,
  IBT1,
  IBT2,
  VSUMESR,
  KBG_N,
  CAPSD,
  CAT0,
  CAT1,
  CAT2,
  CAT3,
  CAT4,
  CAT5,
  ICLR,
  OWL_N,
  ORWD_N,
  OVACC,
  VACC,
  RATR,
  LSD,
  DEL1,
  COMPPAR;
output
  VLENESR_P,
  VST1_P,
  COMPPAR_P,
  BULL5_P,
  END_P,
  PY_P,
  VERR_F,
  PLUTO4_P,
  VSUMESR_P,
  BULL0_P,
  LSD_P,
  STAR2_P,
  SDO,
  PLUTO5_P,
  BULL3_P,
  WATCH_P,
  FBI_P,
  PLUTO2_P,
  MARSSR_P,
  BULL6_P,
  KBG_F,
  STAR0_P,
  PLUTO3_P,
  RATR_P,
  OVACC_P,
  BULL1_P,
  PLUTO0_P,
  STAR3_P,
  VST0_P,
  OWL_F,
  BULL4_P,
  ORWD_F,
  PLUTO1_P,
  ACCRPY_P,
  STAR1_P,
  BULL2_P,
  DEL1_P;
wire
  \[5] ,
  \[45] ,
  \[6] ,
  \[46] ,
  \[7] ,
  \[47] ,
  \[8] ,
  \[48] ,
  \[9] ,
  \[49] ,
  \[20] ,
  \[21] ,
  C1G3,
  \[22] ,
  _1015_m_,
  \[23] ,
  _1214_m_,
  \[24] ,
  \[25] ,
  \[50] ,
  \[26] ,
  \[51] ,
  \[27] ,
  \[28] ,
  \[29] ,
  _254_m__inv,
  \[54] ,
  \[55] ,
  TIMOT,
  \[56] ,
  \[30] ,
  \[31] ,
  C2G5,
  \[32] ,
  \[33] ,
  \[34] ,
  _226_m_,
  \[35] ,
  _873_m_,
  \[36] ,
  \[37] ,
  _44_m__inv,
  \[38] ,
  \[39] ,
  \[10] ,
  \[11] ,
  \[12] ,
  _42_m_,
  _199_m__inv,
  \[13] ,
  \[14] ,
  \[15] ,
  \[40] ,
  \[16] ,
  \[1] ,
  \[41] ,
  \[17] ,
  \[2] ,
  \[42] ,
  \[18] ,
  \[3] ,
  \[43] ,
  \[19] ,
  \[4] ,
  \[44] ;
assign
  \[5]  = (~\[38]  & OWL_N) | (OWL_N & MARSSR),
  \[45]  = \END  & OWL_N,
  \[6]  = (~KBG_N & OWL_N) | (OWL_N & VLENESR),
  \[46]  = C2G5 | ~\[14] ,
  VLENESR_P = \[6] ,
  \[7]  = (\[45]  & VST1) | (OWL_N & VSUMESR),
  \[47]  = ~DEL1 | ~FBI,
  VST1_P = \[25] ,
  COMPPAR_P = \[23] ,
  \[8]  = (\[55]  & \[44] ) | (OWL_N & PLUTO0),
  BULL5_P = \[35] ,
  \[48]  = \[42]  | ~BULL3,
  \[9]  = (\[56]  & \[44] ) | (OWL_N & PLUTO1),
  END_P = \[17] ,
  \[49]  = IBT2 & ~IBT1,
  PY_P = \[16] ,
  VERR_F = \[3] ,
  \[20]  = ~ICLR & VACC,
  \[21]  = (_42_m_ & KBG_N) | ((~_199_m__inv & KBG_N) | ~OWL_N),
  PLUTO4_P = \[12] ,
  C1G3 = (\[50]  & (~IBT0 & ~CAT4)) | ((\[50]  & (IBT0 & ~CAT5)) | ((\[49]  & (~IBT0 & ~CAT2)) | ((\[49]  & (IBT0 & ~CAT3)) | ((\[44]  & (~IBT0 & ~CAT0)) | (\[44]  & (IBT0 & ~CAT1)))))),
  VSUMESR_P = \[7] ,
  \[22]  = ~ICLR & CAPSD,
  _1015_m_ = (\[45]  & \[40] ) | ((\[45]  & VST1) | ((~\[38]  & OWL_N) | (~KBG_N & OWL_N))),
  BULL0_P = \[30] ,
  LSD_P = \[1] ,
  \[23]  = (\[47]  & (COMPPAR & OWL_N)) | (\[41]  & (~COMPPAR & DEL1)),
  _1214_m_ = (\[51]  & OWL_N) | \[30] ,
  \[24]  = (VST1 & (FBI & ~ICLR)) | (\[54]  & VST0),
  STAR2_P = \[28] ,
  \[25]  = (FBI & (PY & ~ICLR)) | (\[54]  & VST1),
  \[50]  = IBT2 & IBT1,
  \[26]  = (~_44_m__inv & STAR0) | (~_254_m__inv & ~STAR0),
  SDO = VST0,
  \[51]  = ~BULL1 | ~BULL0,
  \[27]  = (~_254_m__inv & (~STAR1 & STAR0)) | (\[39]  & STAR1),
  PLUTO5_P = \[13] ,
  BULL3_P = \[33] ,
  \[28]  = (\[43]  & STAR2) | (~_254_m__inv & ~C2G5),
  WATCH_P = \[19] ,
  \[29]  = (~\[43]  & (~_254_m__inv & (C2G5 & ~STAR3))) | ((STAR3 & (~STAR2 & OWL_N)) | (\[43]  & STAR3)),
  FBI_P = \[18] ,
  _254_m__inv = (\[14]  & ~FBI) | ((~FBI & ORWD_N) | ~OWL_N),
  PLUTO2_P = \[10] ,
  \[54]  = ~FBI & ~ICLR,
  \[55]  = _1015_m_ & ~IBT0,
  MARSSR_P = \[5] ,
  TIMOT = ~BULL2 & (BULL1 & (BULL6 & (~BULL5 & (BULL4 & (~BULL3 & ~BULL0))))),
  \[56]  = _1015_m_ & IBT0,
  BULL6_P = \[36] ,
  KBG_F = \[21] ,
  STAR0_P = \[26] ,
  \[30]  = (~BULL0 & (WATCH & OWL_N)) | (BULL0 & (~WATCH & OWL_N)),
  \[31]  = (_1214_m_ & (~\[30]  & BULL0)) | (_1214_m_ & BULL1),
  PLUTO3_P = \[11] ,
  RATR_P = \[4] ,
  C2G5 = STAR2 | (~STAR1 | ~STAR0),
  OVACC_P = \[20] ,
  \[32]  = (_226_m_ & (~_1214_m_ & OWL_N)) | (_1214_m_ & BULL2),
  BULL1_P = \[31] ,
  \[33]  = (~_226_m_ & (~BULL3 & OWL_N)) | (_226_m_ & (BULL3 & OWL_N)),
  PLUTO0_P = \[8] ,
  \[34]  = (~_873_m_ & (BULL4 & OWL_N)) | (_873_m_ & ~BULL4),
  _226_m_ = \[51]  | (~BULL2 | ~WATCH),
  STAR3_P = \[29] ,
  \[35]  = (~_873_m_ & (BULL5 & OWL_N)) | ((_873_m_ & (~\[34]  & ~BULL5)) | (\[34]  & BULL5)),
  _873_m_ = ~_226_m_ & (BULL3 & OWL_N),
  \[36]  = (~\[48]  & (_873_m_ & ~BULL6)) | ((\[48]  & (BULL6 & OWL_N)) | (~_873_m_ & (BULL6 & OWL_N))),
  \[37]  = C2G5 | ~STAR3,
  VST0_P = \[24] ,
  OWL_F = \[15] ,
  _44_m__inv = ~_254_m__inv | ~OWL_N,
  BULL4_P = \[34] ,
  \[38]  = ~TIMOT | ~WATCH,
  ORWD_F = \[14] ,
  \[39]  = (~STAR0 & OWL_N) | ~_44_m__inv,
  PLUTO1_P = \[9] ,
  \[10]  = (\[55]  & \[49] ) | (OWL_N & PLUTO2),
  ACCRPY_P = \[2] ,
  \[11]  = (\[56]  & \[49] ) | (OWL_N & PLUTO3),
  \[12]  = (\[55]  & \[50] ) | (OWL_N & PLUTO4),
  _42_m_ = \[37]  & ~\[14] ,
  _199_m__inv = \[46]  & \[41] ,
  \[13]  = (\[56]  & \[50] ) | (OWL_N & PLUTO5),
  \[14]  = ~C1G3 | ~WATCH,
  STAR1_P = \[27] ,
  \[15]  = \[38]  & (KBG_N & (~\END  & ~ICLR)),
  \[40]  = (~VST0 & ~MMERR) | ~COMPPAR,
  \[16]  = (\[54]  & PY) | (~\[47]  & ~ICLR),
  \[1]  = (~\[41]  & (OWL_N & LSD)) | ((\[41]  & (_42_m_ & ~C2G5)) | (\[37]  & (OWL_N & LSD))),
  \[41]  = FBI & OWL_N,
  \[17]  = (\[41]  & ~_199_m__inv) | \[45] ,
  \[2]  = (\[41]  & ~_199_m__inv) | (OWL_N & ACCRPY),
  \[42]  = ~BULL5 | ~BULL4,
  BULL2_P = \[32] ,
  \[18]  = \[46]  & ~_254_m__inv,
  DEL1_P = \[22] ,
  \[3]  = (\[38]  & (~_199_m__inv & VERR_N)) | ((~TIMOT & (_42_m_ & VERR_N)) | ~OWL_N),
  \[43]  = (~STAR1 & OWL_N) | \[39] ,
  \[19]  = (OVACC & (OWL_N & ~VACC)) | (WATCH & OWL_N),
  \[4]  = (\[45]  & \[40] ) | (OWL_N & RATR),
  \[44]  = ~IBT2 & IBT1;
endmodule

