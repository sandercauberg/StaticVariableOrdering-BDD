module alu4_cl(a, b, c, d, e, f, g, h, i, j, k, l, m, n, o, p, q, r, s, t, u, v);
input
  a,
  b,
  c,
  d,
  e,
  f,
  g,
  h,
  i,
  j,
  k,
  l,
  m,
  n;
output
  o,
  p,
  q,
  r,
  s,
  t,
  u,
  v;
wire
  \[5] ,
  \[99] ,
  \[45] ,
  \[6] ,
  \[46] ,
  \[7] ,
  \[71] ,
  \[47] ,
  \[8] ,
  \[72] ,
  \[48] ,
  \[9] ,
  \[73] ,
  \[49] ,
  \[74] ,
  \[20] ,
  \[75] ,
  \[21] ,
  \[76] ,
  \[22] ,
  \[77] ,
  \[23] ,
  \[78] ,
  \[24] ,
  \[79] ,
  \[25] ,
  \[50] ,
  \[26] ,
  \[27] ,
  \[52] ,
  \[28] ,
  \[53] ,
  \[29] ,
  \[54] ,
  a1,
  a2,
  a3,
  \[55] ,
  b2,
  b3,
  b4,
  \[80] ,
  \[56] ,
  c1,
  c2,
  c4,
  \[57] ,
  d4,
  \[58] ,
  e1,
  e4,
  \[59] ,
  f1,
  g1,
  \[30] ,
  g2,
  g3,
  g4,
  h1,
  \[31] ,
  \[86] ,
  i1,
  \[32] ,
  i3,
  j1,
  \[33] ,
  j4,
  \[34] ,
  k3,
  k4,
  \[35] ,
  l2,
  \[60] ,
  m1,
  \[36] ,
  m2,
  \[61] ,
  \[37] ,
  n3,
  \[62] ,
  \[38] ,
  o3,
  p0,
  \[63] ,
  p1,
  \[39] ,
  p2,
  q0,
  \[64] ,
  q2,
  \[10] ,
  q3,
  \[65] ,
  r1,
  \[11] ,
  r3,
  s1,
  \[12] ,
  s3,
  t0,
  \[67] ,
  \[13] ,
  \[68] ,
  u2,
  \[14] ,
  u3,
  v0,
  \[69] ,
  v2,
  \[15] ,
  \[0] ,
  \[94] ,
  w0,
  w1,
  \[40] ,
  w2,
  \[16] ,
  w3,
  \[1] ,
  \[41] ,
  \[17] ,
  x3,
  \[2] ,
  \[96] ,
  y0,
  y1,
  \[42] ,
  y2,
  \[18] ,
  \[3] ,
  \[97] ,
  z0,
  \[43] ,
  z2,
  z3,
  \[4] ,
  \[98] ,
  \[44] ;
assign
  \[5]  = h & d,
  \[99]  = w0 & ~n,
  \[45]  = v0 & n,
  \[6]  = (~\[44]  & (~\[11]  & (~v0 & (~p0 & (~r1 & n))))) | ((\[97]  & (~\[60]  & (\[44]  & ~r1))) | ((\[60]  & (~p0 & (r1 & n))) | ((~\[9]  & (t0 & (~h1 & d))) | ((\[11]  & (~p0 & ~\[4] )) | ((\[11]  & (~s1 & \[5] )) | ((\[9]  & (c1 & d)) | ((~\[50]  & p0) | ((\[21]  & v0) | i1)))))))),
  \[46]  = ~n & l,
  \[7]  = (~\[22]  & (\[20]  & (\[8]  & \[4] ))) | (\[20]  & (\[8]  & (a2 & \[4] ))),
  \[71]  = \[12]  & r1,
  \[47]  = z0 | t0,
  \[8]  = (~n3 & ~a) | k3,
  \[72]  = 0,
  \[48]  = (b4 & ~j) | k4,
  \[9]  = g2 & n,
  \[73]  = r1 & (~n & k),
  \[49]  = \[17]  | v2,
  \[74]  = c4 & ~k,
  \[20]  = q2 | p2,
  \[75]  = ~m2 & ~i3,
  o = \[0] ,
  \[21]  = (y0 & (r1 & (n & ~d))) | (~\[49]  & (b4 & ~t0)),
  p = \[1] ,
  q = \[2] ,
  r = \[3] ,
  s = \[4] ,
  t = \[5] ,
  u = \[6] ,
  v = \[7] ,
  \[76]  = h1 & d,
  \[22]  = g | c,
  \[77]  = 0,
  \[23]  = (u2 & v2) | ~\[86] ,
  \[78]  = \[27]  & p1,
  \[24]  = j & ~i,
  \[79]  = \[45]  & r1,
  \[25]  = ~w3 | ~i3,
  \[50]  = \[26]  | ~w1,
  \[26]  = \[15]  | ~l2,
  \[27]  = ~n & j,
  \[52]  = \[12]  & l,
  \[28]  = m2 | b,
  \[53]  = \[27]  & (u3 & s1),
  \[29]  = (z0 & h1) | ~\[60] ,
  \[54]  = u3 & q0,
  a1 = (\[86]  & w2) | (u2 & v2),
  a2 = g & c,
  a3 = (~v2 & x3) | (v2 & ~x3),
  \[55]  = n & ~l,
  b2 = c2 & ~m1,
  b3 = (\[58]  & \[28] ) | \[69] ,
  b4 = u3 & n,
  \[80]  = \[12]  & s1,
  \[56]  = ~s1 & ~j,
  c1 = (\[35]  & b3) | \[67] ,
  c2 = (q0 & (l & ~k)) | (\[24]  & ~l),
  c4 = \[33]  & j,
  \[57]  = b2 & n,
  d4 = (\[52]  & (k & i)) | ((\[40]  & ~u3) | \[54] ),
  \[58]  = i3 & a,
  e1 = (\[22]  & \[14] ) | a2,
  e4 = (\[56]  & (n & k)) | (\[99]  & s1),
  \[59]  = t0 | d,
  f1 = ~j & ~i,
  g1 = (~a3 & x3) | (a3 & c),
  \[30]  = \[76]  | ~\[39] ,
  g2 = (~q0 & (k & l)) | (f1 & l),
  g3 = (~\[38]  & (~\[9]  & (q3 & i3))) | ((\[11]  & (~k3 & a)) | ((\[9]  & (~i3 & a)) | ((\[9]  & (i3 & ~a)) | ((\[96]  & i3) | ((\[96]  & a) | ((\[79]  & ~a) | ((\[57]  & ~i3) | ((\[38]  & ~q3) | ((\[13]  & ~q3) | ((\[13]  & ~a) | ((\[11]  & n3) | (z3 & ~i3)))))))))))),
  g4 = (~g & c) | ((~g & ~j4) | (c & ~j4)),
  h1 = (~k4 & (f1 & (s1 & (n & c)))) | ((~g4 & (b4 & (b2 & \[4] ))) | ((g4 & (b4 & (b2 & ~\[4] ))) | ((\[61]  & (\[41]  & ~d)) | ((k4 & \[5] ) | ((e4 & \[5] ) | ((e4 & ~\[4] ) | (d4 & ~h))))))),
  \[31]  = (t0 & d) | ~\[59] ,
  \[86]  = u2 | v2,
  i1 = (y2 & u2) | z2,
  \[32]  = \[16]  | m2,
  i3 = (\[40]  & (~\[8]  & ~d4)) | ((\[94]  & ~a) | ((~\[8]  & e4) | ((k4 & k3) | ((e4 & a) | (d4 & ~e))))),
  j1 = (\[55]  & (q0 & ~k)) | (\[12]  & (p1 & k)),
  \[33]  = p1 & n,
  j4 = (\[62]  & n3) | \[98] ,
  \[34]  = s3,
  k3 = e & a,
  k4 = (\[57]  & q0) | ((\[9]  & ~k) | (u3 & f1)),
  \[35]  = y1 | c,
  l2 = (~\[38]  & (\[28]  & (\[16]  & (\[10]  & (~\[9]  & (~q2 & ~k3)))))) | ((~\[57]  & (\[55]  & (~\[43]  & (~o3 & b)))) | ((~\[55]  & (\[20]  & (\[11]  & k3))) | ((\[79]  & (\[28]  & a)) | ((\[69]  & (\[58]  & \[9] )) | ((\[58]  & (~\[28]  & \[9] )) | ((\[55]  & (~\[20]  & \[11] )) | ((\[44]  & (\[16]  & m2)) | ((\[28]  & (\[9]  & ~b3)) | ((~\[20]  & (\[11]  & ~k3)) | ((\[79]  & ~\[36] ) | ((\[75]  & \[57] ) | ((\[75]  & ~\[37] ) | ((\[43]  & ~z2) | ((\[38]  & ~\[17] ) | (\[13]  & ~x3))))))))))))))),
  \[60]  = z0 | h1,
  m1 = ~k & ~i,
  \[36]  = b | a,
  m2 = (~\[40]  & (\[33]  & (~m1 & a))) | ((\[40]  & (~\[20]  & (~d4 & ~n3))) | ((\[40]  & (\[20]  & (j4 & ~d4))) | ((\[94]  & ~b) | ((\[48]  & q2) | ((e4 & ~p2) | (d4 & ~f)))))),
  \[61]  = c2 | f1,
  \[37]  = ~w3 | ~q3,
  n3 = e & ~a,
  \[62]  = f | ~b,
  \[38]  = b4 & v0,
  o3 = (~\[63]  & ~r3) | (\[63]  & r3),
  p0 = (~\[38]  & (~\[29]  & (~\[18]  & (~\[9]  & (~i1 & ~a1))))) | ((~\[96]  & (\[11]  & (e1 & \[4] ))) | ((\[97]  & (\[57]  & \[29] )) | ((\[96]  & (\[11]  & ~\[4] )) | ((\[79]  & (~\[31]  & ~y0)) | ((\[57]  & (~\[29]  & y1)) | ((\[49]  & (\[38]  & ~\[18] )) | ((\[44]  & (\[32]  & ~\[29] )) | ((~\[31]  & (\[13]  & ~g1)) | ((~\[30]  & (\[13]  & g1)) | ((~\[30]  & (\[9]  & ~c1)) | ((\[30]  & (\[9]  & c1)) | ((\[11]  & (~e1 & ~\[4] )) | ((\[96]  & ~\[31] ) | ((\[29]  & i1) | ((\[21]  & v0) | (\[18]  & a1)))))))))))))))),
  \[63]  = ~q3 | ~a,
  p1 = l & ~i,
  \[39]  = h1 | d,
  p2 = ~f & ~b,
  q0 = j & i,
  \[64]  = b4 & q0,
  q2 = f & b,
  \[10]  = (~s3 & r3) | (s3 & ~r3),
  q3 = (\[64]  & \[58] ) | ((\[13]  & ~i3) | ((z3 & k3) | ((c4 & i3) | (c4 & a)))),
  \[65]  = \[46]  & ~w0,
  r1 = (l & k) | m1,
  \[11]  = w0 & n,
  r3 = (\[69]  & \[64] ) | ((\[28]  & c4) | ((\[13]  & ~m2) | (z3 & q2))),
  s1 = (~l & (~k & i)) | (k & ~i),
  \[12]  = ~n & ~j,
  s3 = (\[74]  & q2) | (~r3 & z3),
  t0 = (\[76]  & \[64] ) | ((\[39]  & c4) | ((\[13]  & ~h1) | (z3 & \[5] ))),
  \[67]  = y1 & c,
  \[13]  = b4 & f1,
  \[68]  = \[56]  & (u3 & ~e4),
  u2 = (\[74]  & a2) | (z3 & ~v2),
  \[14]  = (~p2 & k3) | q2,
  u3 = ~l & k,
  v0 = q0 & k,
  \[69]  = m2 & b,
  v2 = (\[67]  & \[64] ) | ((\[35]  & c4) | ((\[13]  & ~y1) | (z3 & a2))),
  \[15]  = ~g3 | m,
  \[0]  = (~\[99]  & (~\[8]  & (i3 & ~n))) | ((~\[73]  & (\[52]  & ~\[8] )) | ((~g3 & (n & ~m)) | ((\[80]  & ~i3) | ((\[78]  & n3) | ((\[73]  & a) | ((\[71]  & i3) | ((\[68]  & ~e) | ((\[65]  & k3) | ((\[53]  & \[8] ) | ((g3 & m) | j1)))))))))),
  \[94]  = (\[52]  & \[41] ) | (\[41]  & ~l),
  w0 = ~k & (~j & i),
  w1 = (~\[45]  & (~\[23]  & (~\[9]  & (~y2 & (~z2 & ~w2))))) | ((\[97]  & (\[45]  & (\[36]  & c))) | ((~\[96]  & (~\[22]  & (\[14]  & \[11] ))) | ((\[96]  & (\[11]  & e1)) | ((\[67]  & (\[45]  & \[17] )) | ((\[67]  & (\[9]  & b3)) | ((\[61]  & (~\[35]  & a3)) | ((\[44]  & (\[32]  & ~y2)) | ((~\[35]  & (\[9]  & b3)) | ((\[35]  & (\[9]  & ~c1)) | ((\[22]  & (\[11]  & ~e1)) | ((\[14]  & (\[11]  & a2)) | ((\[13]  & (~a3 & c)) | ((\[97]  & \[57] ) | ((\[96]  & \[35] ) | ((~\[49]  & \[38] ) | ((\[45]  & y0) | ((\[23]  & w2) | (y2 & z2)))))))))))))))))),
  \[40]  = \[24]  & n,
  w2 = (~\[37]  & r3) | (s3 & r3),
  \[16]  = i3 | m1,
  w3 = (\[74]  & k3) | (~q3 & z3),
  \[1]  = (~\[99]  & (~\[20]  & (m2 & ~n))) | ((~\[73]  & (\[52]  & ~\[20] )) | ((\[98]  & \[78] ) | ((\[80]  & ~m2) | ((\[73]  & b) | ((\[71]  & m2) | ((\[68]  & ~f) | ((\[65]  & q2) | ((\[53]  & \[20] ) | ((~\[15]  & ~l2) | ((\[15]  & l2) | j1)))))))))),
  \[41]  = m1 & ~n,
  \[17]  = r3 | q3,
  x3 = (~\[63]  & ~o3) | (o3 & b),
  \[2]  = (~\[80]  & (\[22]  & (y1 & ~n))) | ((~\[73]  & (\[52]  & (\[22]  & ~a2))) | ((\[80]  & ~y1) | ((\[78]  & g) | ((\[73]  & c) | ((\[71]  & ~\[22] ) | ((\[68]  & ~g) | ((\[65]  & a2) | ((\[53]  & ~\[22] ) | ((\[53]  & a2) | ((~\[26]  & ~w1) | ((\[26]  & w1) | j1))))))))))),
  \[96]  = \[55]  & (~u3 & ~q0),
  y0 = ~\[36]  & ~c,
  y1 = (\[40]  & (\[22]  & (~j4 & (~d4 & ~a2)))) | ((~\[40]  & (\[33]  & (~m1 & b))) | ((\[40]  & (~g4 & (~d4 & a2))) | ((\[40]  & (~\[22]  & ~g4)) | ((\[94]  & ~c) | ((\[48]  & a2) | ((\[22]  & e4) | (d4 & ~g))))))),
  \[42]  = 0,
  y2 = (~y1 & ~u2) | (y1 & u2),
  \[18]  = (z0 & t0) | ~\[47] ,
  \[3]  = (~\[80]  & (h1 & (~\[4]  & ~n))) | ((~\[73]  & (\[52]  & ~\[4] )) | ((\[80]  & ~h1) | ((\[78]  & h) | ((\[73]  & d) | ((\[71]  & h1) | ((\[68]  & ~h) | ((\[65]  & \[5] ) | ((\[53]  & \[4] ) | ((~\[50]  & ~p0) | ((\[50]  & p0) | j1)))))))))),
  \[97]  = \[75]  & ~y1,
  z0 = (\[74]  & \[5] ) | (z3 & ~t0),
  \[43]  = u3 & e4,
  z2 = (\[34]  & m2) | ~\[25] ,
  z3 = b4 & (~j & i),
  \[4]  = (~h & ~d) | \[5] ,
  \[98]  = f & ~b,
  \[44]  = c2 & n;
endmodule

